-- this file was generated with hex2rom written by daniel wallner

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
	port(
		ce_n	: in std_logic;
		oe_n	: in std_logic;
		a	: in std_logic_vector(13 downto 0);
		d	: out std_logic_vector(7 downto 0)
	);
end rom;

architecture rtl of rom is
	subtype rom_word is std_logic_vector(7 downto 0);
	type rom_table is array(0 to 16383) of rom_word;
	constant rom: rom_table := rom_table'(
		"01011111",	-- 0x0000
		"01011111",	-- 0x0001
		"01011111",	-- 0x0002
		"01000000",	-- 0x0003
		"11111110",	-- 0x0004
		"00000000",	-- 0x0005
		"00000010",	-- 0x0006
		"00000000",	-- 0x0007
		"00010000",	-- 0x0008
		"00000000",	-- 0x0009
		"00000000",	-- 0x000a
		"00001010",	-- 0x000b
		"00101011",	-- 0x000c
		"00100111",	-- 0x000d
		"00011110",	-- 0x000e
		"00011000",	-- 0x000f
		"00010110",	-- 0x0010
		"00010010",	-- 0x0011
		"00010010",	-- 0x0012
		"00001111",	-- 0x0013
		"00001110",	-- 0x0014
		"00001110",	-- 0x0015
		"00001101",	-- 0x0016
		"00001100",	-- 0x0017
		"00001100",	-- 0x0018
		"00001100",	-- 0x0019
		"00001100",	-- 0x001a
		"00001100",	-- 0x001b
		"00001100",	-- 0x001c
		"01001100",	-- 0x001d
		"01001001",	-- 0x001e
		"01000101",	-- 0x001f
		"00111010",	-- 0x0020
		"00101111",	-- 0x0021
		"00100111",	-- 0x0022
		"00100001",	-- 0x0023
		"00011010",	-- 0x0024
		"00010110",	-- 0x0025
		"00010110",	-- 0x0026
		"00010101",	-- 0x0027
		"00010010",	-- 0x0028
		"00010010",	-- 0x0029
		"00010010",	-- 0x002a
		"00010010",	-- 0x002b
		"00010010",	-- 0x002c
		"00010010",	-- 0x002d
		"01011011",	-- 0x002e
		"01011000",	-- 0x002f
		"01011000",	-- 0x0030
		"01010000",	-- 0x0031
		"01001010",	-- 0x0032
		"01000000",	-- 0x0033
		"00110101",	-- 0x0034
		"00101101",	-- 0x0035
		"00100111",	-- 0x0036
		"00100101",	-- 0x0037
		"00100010",	-- 0x0038
		"00011101",	-- 0x0039
		"00011101",	-- 0x003a
		"00011101",	-- 0x003b
		"00011101",	-- 0x003c
		"00011101",	-- 0x003d
		"00011101",	-- 0x003e
		"01011101",	-- 0x003f
		"01011100",	-- 0x0040
		"01011011",	-- 0x0041
		"01011000",	-- 0x0042
		"01010110",	-- 0x0043
		"01001110",	-- 0x0044
		"01000111",	-- 0x0045
		"00111111",	-- 0x0046
		"00111000",	-- 0x0047
		"00110101",	-- 0x0048
		"00110001",	-- 0x0049
		"00101010",	-- 0x004a
		"00101010",	-- 0x004b
		"00101010",	-- 0x004c
		"00101010",	-- 0x004d
		"00101010",	-- 0x004e
		"00101010",	-- 0x004f
		"01011110",	-- 0x0050
		"01011110",	-- 0x0051
		"01011110",	-- 0x0052
		"01011100",	-- 0x0053
		"01011011",	-- 0x0054
		"01010111",	-- 0x0055
		"01010010",	-- 0x0056
		"01001100",	-- 0x0057
		"01000110",	-- 0x0058
		"01000011",	-- 0x0059
		"00111110",	-- 0x005a
		"00111000",	-- 0x005b
		"00111000",	-- 0x005c
		"00111000",	-- 0x005d
		"00111000",	-- 0x005e
		"00111000",	-- 0x005f
		"00111000",	-- 0x0060
		"01011110",	-- 0x0061
		"01011110",	-- 0x0062
		"01011111",	-- 0x0063
		"01011110",	-- 0x0064
		"01011110",	-- 0x0065
		"01011010",	-- 0x0066
		"01010111",	-- 0x0067
		"01010011",	-- 0x0068
		"01001111",	-- 0x0069
		"01001011",	-- 0x006a
		"01001001",	-- 0x006b
		"01000011",	-- 0x006c
		"01000011",	-- 0x006d
		"01000011",	-- 0x006e
		"01000011",	-- 0x006f
		"01000011",	-- 0x0070
		"01000011",	-- 0x0071
		"01100000",	-- 0x0072
		"01100000",	-- 0x0073
		"01100000",	-- 0x0074
		"01100000",	-- 0x0075
		"01011111",	-- 0x0076
		"01011110",	-- 0x0077
		"01011101",	-- 0x0078
		"01011011",	-- 0x0079
		"01011010",	-- 0x007a
		"01011000",	-- 0x007b
		"01010110",	-- 0x007c
		"01010011",	-- 0x007d
		"01010011",	-- 0x007e
		"01010011",	-- 0x007f
		"01010011",	-- 0x0080
		"01010011",	-- 0x0081
		"01010011",	-- 0x0082
		"01100001",	-- 0x0083
		"01100000",	-- 0x0084
		"01100000",	-- 0x0085
		"01100000",	-- 0x0086
		"01100000",	-- 0x0087
		"01100000",	-- 0x0088
		"01011111",	-- 0x0089
		"01011110",	-- 0x008a
		"01011110",	-- 0x008b
		"01011101",	-- 0x008c
		"01011100",	-- 0x008d
		"01011011",	-- 0x008e
		"01011011",	-- 0x008f
		"01011011",	-- 0x0090
		"01011011",	-- 0x0091
		"01011011",	-- 0x0092
		"01011011",	-- 0x0093
		"01100001",	-- 0x0094
		"01100001",	-- 0x0095
		"01100001",	-- 0x0096
		"01100001",	-- 0x0097
		"01100001",	-- 0x0098
		"01100001",	-- 0x0099
		"01100000",	-- 0x009a
		"01011111",	-- 0x009b
		"01011111",	-- 0x009c
		"01011111",	-- 0x009d
		"01011111",	-- 0x009e
		"01011110",	-- 0x009f
		"01011110",	-- 0x00a0
		"01011110",	-- 0x00a1
		"01011110",	-- 0x00a2
		"01011110",	-- 0x00a3
		"01011110",	-- 0x00a4
		"01100001",	-- 0x00a5
		"01100001",	-- 0x00a6
		"01100001",	-- 0x00a7
		"01100001",	-- 0x00a8
		"01100001",	-- 0x00a9
		"01100001",	-- 0x00aa
		"01100001",	-- 0x00ab
		"01100001",	-- 0x00ac
		"01100001",	-- 0x00ad
		"01100000",	-- 0x00ae
		"01100001",	-- 0x00af
		"01100001",	-- 0x00b0
		"01100001",	-- 0x00b1
		"01100001",	-- 0x00b2
		"01100001",	-- 0x00b3
		"01100001",	-- 0x00b4
		"01100001",	-- 0x00b5
		"01100001",	-- 0x00b6
		"01100001",	-- 0x00b7
		"01100001",	-- 0x00b8
		"01100001",	-- 0x00b9
		"01100001",	-- 0x00ba
		"01100001",	-- 0x00bb
		"01100001",	-- 0x00bc
		"01100001",	-- 0x00bd
		"01100001",	-- 0x00be
		"01100001",	-- 0x00bf
		"01100001",	-- 0x00c0
		"01100001",	-- 0x00c1
		"01100001",	-- 0x00c2
		"01100001",	-- 0x00c3
		"01100001",	-- 0x00c4
		"01100001",	-- 0x00c5
		"01100001",	-- 0x00c6
		"00000000",	-- 0x00c7
		"10000000",	-- 0x00c8
		"00000010",	-- 0x00c9
		"00000010",	-- 0x00ca
		"00100101",	-- 0x00cb
		"00001010",	-- 0x00cc
		"00000011",	-- 0x00cd
		"00010001",	-- 0x00ce
		"00011010",	-- 0x00cf
		"00000100",	-- 0x00d0
		"00010011",	-- 0x00d1
		"00011111",	-- 0x00d2
		"00000100",	-- 0x00d3
		"00010100",	-- 0x00d4
		"00100110",	-- 0x00d5
		"00000101",	-- 0x00d6
		"00010101",	-- 0x00d7
		"00101000",	-- 0x00d8
		"00000101",	-- 0x00d9
		"00010110",	-- 0x00da
		"00101011",	-- 0x00db
		"00000110",	-- 0x00dc
		"00010111",	-- 0x00dd
		"00101110",	-- 0x00de
		"00000110",	-- 0x00df
		"00011001",	-- 0x00e0
		"00110000",	-- 0x00e1
		"00001010",	-- 0x00e2
		"00100010",	-- 0x00e3
		"00110010",	-- 0x00e4
		"00001101",	-- 0x00e5
		"00100000",	-- 0x00e6
		"00110101",	-- 0x00e7
		"00001111",	-- 0x00e8
		"00100110",	-- 0x00e9
		"00111101",	-- 0x00ea
		"00110000",	-- 0x00eb
		"00111110",	-- 0x00ec
		"01001100",	-- 0x00ed
		"00000010",	-- 0x00ee
		"10000000",	-- 0x00ef
		"00000101",	-- 0x00f0
		"00000001",	-- 0x00f1
		"00000000",	-- 0x00f2
		"00000100",	-- 0x00f3
		"10000000",	-- 0x00f4
		"10000000",	-- 0x00f5
		"01011010",	-- 0x00f6
		"01011010",	-- 0x00f7
		"01011010",	-- 0x00f8
		"01011010",	-- 0x00f9
		"10000000",	-- 0x00fa
		"10000000",	-- 0x00fb
		"01001101",	-- 0x00fc
		"01001101",	-- 0x00fd
		"01001101",	-- 0x00fe
		"01001101",	-- 0x00ff
		"10000000",	-- 0x0100
		"10000000",	-- 0x0101
		"00110011",	-- 0x0102
		"00110011",	-- 0x0103
		"00110011",	-- 0x0104
		"00110011",	-- 0x0105
		"10000000",	-- 0x0106
		"10000000",	-- 0x0107
		"00110011",	-- 0x0108
		"00110011",	-- 0x0109
		"00110011",	-- 0x010a
		"00110011",	-- 0x010b
		"10000000",	-- 0x010c
		"10000000",	-- 0x010d
		"00110011",	-- 0x010e
		"00110011",	-- 0x010f
		"00110011",	-- 0x0110
		"00110011",	-- 0x0111
		"00011000",	-- 0x0112
		"00010000",	-- 0x0113
		"01100111",	-- 0x0114
		"00100000",	-- 0x0115
		"01011100",	-- 0x0116
		"00101111",	-- 0x0117
		"01001011",	-- 0x0118
		"00111111",	-- 0x0119
		"00111011",	-- 0x011a
		"01001110",	-- 0x011b
		"00110101",	-- 0x011c
		"01011110",	-- 0x011d
		"00101001",	-- 0x011e
		"01101101",	-- 0x011f
		"00011110",	-- 0x0120
		"01111101",	-- 0x0121
		"00010111",	-- 0x0122
		"10001101",	-- 0x0123
		"00001111",	-- 0x0124
		"10011101",	-- 0x0125
		"00001110",	-- 0x0126
		"10101101",	-- 0x0127
		"00001101",	-- 0x0128
		"10111101",	-- 0x0129
		"00001010",	-- 0x012a
		"11001101",	-- 0x012b
		"00001001",	-- 0x012c
		"00000010",	-- 0x012d
		"10000000",	-- 0x012e
		"00000110",	-- 0x012f
		"11111111",	-- 0x0130
		"10010010",	-- 0x0131
		"01110010",	-- 0x0132
		"01011101",	-- 0x0133
		"01001111",	-- 0x0134
		"01000100",	-- 0x0135
		"00111100",	-- 0x0136
		"10011100",	-- 0x0137
		"01000000",	-- 0x0138
		"11111111",	-- 0x0139
		"10100000",	-- 0x013a
		"01000000",	-- 0x013b
		"01000110",	-- 0x013c
		"00010000",	-- 0x013d
		"10101001",	-- 0x013e
		"10010100",	-- 0x013f
		"01010011",	-- 0x0140
		"10000000",	-- 0x0141
		"10101001",	-- 0x0142
		"01001110",	-- 0x0143
		"00101010",	-- 0x0144
		"00011110",	-- 0x0145
		"00010001",	-- 0x0146
		"00100110",	-- 0x0147
		"11000000",	-- 0x0148
		"01100000",	-- 0x0149
		"01010000",	-- 0x014a
		"01000100",	-- 0x014b
		"00101010",	-- 0x014c
		"01100000",	-- 0x014d
		"10000000",	-- 0x014e
		"00001111",	-- 0x014f
		"00000110",	-- 0x0150
		"00000110",	-- 0x0151
		"00000110",	-- 0x0152
		"00000110",	-- 0x0153
		"00000001",	-- 0x0154
		"00010011",	-- 0x0155
		"00001011",	-- 0x0156
		"00000000",	-- 0x0157
		"00000111",	-- 0x0158
		"00001001",	-- 0x0159
		"00010011",	-- 0x015a
		"00011001",	-- 0x015b
		"00100000",	-- 0x015c
		"00100101",	-- 0x015d
		"00101011",	-- 0x015e
		"00111011",	-- 0x015f
		"01001110",	-- 0x0160
		"01101001",	-- 0x0161
		"10000000",	-- 0x0162
		"00000001",	-- 0x0163
		"00000000",	-- 0x0164
		"00000001",	-- 0x0165
		"00011010",	-- 0x0166
		"10000000",	-- 0x0167
		"00000000",	-- 0x0168
		"10000000",	-- 0x0169
		"00000110",	-- 0x016a
		"01000111",	-- 0x016b
		"01000111",	-- 0x016c
		"01001001",	-- 0x016d
		"01010110",	-- 0x016e
		"00110000",	-- 0x016f
		"00110000",	-- 0x0170
		"00110000",	-- 0x0171
		"00000000",	-- 0x0172
		"10000000",	-- 0x0173
		"00000110",	-- 0x0174
		"01000010",	-- 0x0175
		"01000010",	-- 0x0176
		"01010111",	-- 0x0177
		"01000011",	-- 0x0178
		"01000101",	-- 0x0179
		"01000101",	-- 0x017a
		"01000101",	-- 0x017b
		"00011111",	-- 0x017c
		"11000000",	-- 0x017d
		"00110000",	-- 0x017e
		"00110000",	-- 0x017f
		"01100100",	-- 0x0180
		"00111111",	-- 0x0181
		"00100000",	-- 0x0182
		"00000110",	-- 0x0183
		"00000000",	-- 0x0184
		"00011111",	-- 0x0185
		"11000000",	-- 0x0186
		"00000000",	-- 0x0187
		"00000000",	-- 0x0188
		"00000000",	-- 0x0189
		"00000000",	-- 0x018a
		"00000000",	-- 0x018b
		"00000000",	-- 0x018c
		"00000000",	-- 0x018d
		"00001110",	-- 0x018e
		"00011111",	-- 0x018f
		"10000000",	-- 0x0190
		"00111110",	-- 0x0191
		"10000000",	-- 0x0192
		"01011101",	-- 0x0193
		"01100000",	-- 0x0194
		"01111100",	-- 0x0195
		"01000000",	-- 0x0196
		"10011100",	-- 0x0197
		"00101000",	-- 0x0198
		"10111100",	-- 0x0199
		"00010100",	-- 0x019a
		"11011100",	-- 0x019b
		"00000110",	-- 0x019c
		"11101000",	-- 0x019d
		"00000000",	-- 0x019e
		"00001110",	-- 0x019f
		"00011111",	-- 0x01a0
		"01101100",	-- 0x01a1
		"00111110",	-- 0x01a2
		"01101010",	-- 0x01a3
		"01011101",	-- 0x01a4
		"01010100",	-- 0x01a5
		"01111100",	-- 0x01a6
		"01001000",	-- 0x01a7
		"10011100",	-- 0x01a8
		"00011100",	-- 0x01a9
		"10111100",	-- 0x01aa
		"00010010",	-- 0x01ab
		"11011100",	-- 0x01ac
		"00000111",	-- 0x01ad
		"11101000",	-- 0x01ae
		"00000000",	-- 0x01af
		"00001110",	-- 0x01b0
		"00011111",	-- 0x01b1
		"00000000",	-- 0x01b2
		"00111110",	-- 0x01b3
		"00000000",	-- 0x01b4
		"01011101",	-- 0x01b5
		"00000000",	-- 0x01b6
		"01111100",	-- 0x01b7
		"00000000",	-- 0x01b8
		"10011100",	-- 0x01b9
		"00000000",	-- 0x01ba
		"10111100",	-- 0x01bb
		"00000000",	-- 0x01bc
		"11011100",	-- 0x01bd
		"00000000",	-- 0x01be
		"11101000",	-- 0x01bf
		"00000000",	-- 0x01c0
		"00001110",	-- 0x01c1
		"00011111",	-- 0x01c2
		"00000000",	-- 0x01c3
		"00111110",	-- 0x01c4
		"00000000",	-- 0x01c5
		"01011101",	-- 0x01c6
		"00000000",	-- 0x01c7
		"01111100",	-- 0x01c8
		"00000000",	-- 0x01c9
		"10011100",	-- 0x01ca
		"00000000",	-- 0x01cb
		"10111100",	-- 0x01cc
		"00000000",	-- 0x01cd
		"11011100",	-- 0x01ce
		"00000000",	-- 0x01cf
		"11101000",	-- 0x01d0
		"00000000",	-- 0x01d1
		"00111000",	-- 0x01d2
		"01100000",	-- 0x01d3
		"01111101",	-- 0x01d4
		"01111101",	-- 0x01d5
		"01111101",	-- 0x01d6
		"01111101",	-- 0x01d7
		"00000110",	-- 0x01d8
		"00100110",	-- 0x01d9
		"00000000",	-- 0x01da
		"01010001",	-- 0x01db
		"00000000",	-- 0x01dc
		"10000110",	-- 0x01dd
		"00000000",	-- 0x01de
		"10110011",	-- 0x01df
		"00000000",	-- 0x01e0
		"00011000",	-- 0x01e1
		"01100000",	-- 0x01e2
		"01100110",	-- 0x01e3
		"00101010",	-- 0x01e4
		"00101000",	-- 0x01e5
		"00110011",	-- 0x01e6
		"00111000",	-- 0x01e7
		"01010000",	-- 0x01e8
		"00000010",	-- 0x01e9
		"00000011",	-- 0x01ea
		"00000101",	-- 0x01eb
		"00001001",	-- 0x01ec
		"00001011",	-- 0x01ed
		"00011010",	-- 0x01ee
		"00000010",	-- 0x01ef
		"00000000",	-- 0x01f0
		"00000010",	-- 0x01f1
		"11011010",	-- 0x01f2
		"11011010",	-- 0x01f3
		"11011010",	-- 0x01f4
		"00000010",	-- 0x01f5
		"00000000",	-- 0x01f6
		"00000010",	-- 0x01f7
		"01100010",	-- 0x01f8
		"01100010",	-- 0x01f9
		"01100010",	-- 0x01fa
		"00000010",	-- 0x01fb
		"01010001",	-- 0x01fc
		"00100110",	-- 0x01fd
		"11100100",	-- 0x01fe
		"00100110",	-- 0x01ff
		"00000110",	-- 0x0200
		"00101001",	-- 0x0201
		"01111010",	-- 0x0202
		"01010010",	-- 0x0203
		"01011100",	-- 0x0204
		"01111011",	-- 0x0205
		"00111101",	-- 0x0206
		"10100100",	-- 0x0207
		"00111101",	-- 0x0208
		"00001000",	-- 0x0209
		"00101000",	-- 0x020a
		"01000000",	-- 0x020b
		"00111100",	-- 0x020c
		"01110011",	-- 0x020d
		"01010000",	-- 0x020e
		"01111111",	-- 0x020f
		"01100100",	-- 0x0210
		"01111111",	-- 0x0211
		"01111000",	-- 0x0212
		"01111111",	-- 0x0213
		"00010010",	-- 0x0214
		"00001010",	-- 0x0215
		"11111101",	-- 0x0216
		"00010100",	-- 0x0217
		"11111101",	-- 0x0218
		"00011111",	-- 0x0219
		"11111101",	-- 0x021a
		"00101001",	-- 0x021b
		"11111101",	-- 0x021c
		"00110011",	-- 0x021d
		"00011010",	-- 0x021e
		"00111101",	-- 0x021f
		"00000000",	-- 0x0220
		"01001000",	-- 0x0221
		"00000000",	-- 0x0222
		"01010010",	-- 0x0223
		"00000000",	-- 0x0224
		"01011100",	-- 0x0225
		"00000000",	-- 0x0226
		"01100110",	-- 0x0227
		"00000000",	-- 0x0228
		"00001010",	-- 0x0229
		"00000101",	-- 0x022a
		"00001010",	-- 0x022b
		"00000101",	-- 0x022c
		"00011010",	-- 0x022d
		"00011010",	-- 0x022e
		"00011010",	-- 0x022f
		"00011010",	-- 0x0230
		"00101011",	-- 0x0231
		"00010110",	-- 0x0232
		"00010000",	-- 0x0233
		"01000000",	-- 0x0234
		"01000001",	-- 0x0235
		"01100001",	-- 0x0236
		"10010111",	-- 0x0237
		"00010000",	-- 0x0238
		"01000000",	-- 0x0239
		"01000001",	-- 0x023a
		"01100001",	-- 0x023b
		"01101100",	-- 0x023c
		"00101011",	-- 0x023d
		"00010110",	-- 0x023e
		"00010000",	-- 0x023f
		"01000000",	-- 0x0240
		"01000001",	-- 0x0241
		"01101100",	-- 0x0242
		"10100001",	-- 0x0243
		"00010000",	-- 0x0244
		"01000000",	-- 0x0245
		"01000001",	-- 0x0246
		"01010110",	-- 0x0247
		"01100001",	-- 0x0248
		"00001001",	-- 0x0249
		"00001001",	-- 0x024a
		"00000110",	-- 0x024b
		"00010000",	-- 0x024c
		"00001011",	-- 0x024d
		"11111110",	-- 0x024e
		"11111110",	-- 0x024f
		"11111110",	-- 0x0250
		"11111110",	-- 0x0251
		"11111110",	-- 0x0252
		"01000000",	-- 0x0253
		"01010000",	-- 0x0254
		"01111010",	-- 0x0255
		"01111010",	-- 0x0256
		"01111010",	-- 0x0257
		"00110001",	-- 0x0258
		"00110001",	-- 0x0259
		"00110001",	-- 0x025a
		"00000000",	-- 0x025b
		"00000000",	-- 0x025c
		"00000000",	-- 0x025d
		"00000000",	-- 0x025e
		"00001000",	-- 0x025f
		"00000000",	-- 0x0260
		"00000000",	-- 0x0261
		"00000000",	-- 0x0262
		"00001101",	-- 0x0263
		"00001101",	-- 0x0264
		"00001101",	-- 0x0265
		"00001101",	-- 0x0266
		"00001000",	-- 0x0267
		"10000000",	-- 0x0268
		"11111111",	-- 0x0269
		"10011010",	-- 0x026a
		"11010111",	-- 0x026b
		"10110011",	-- 0x026c
		"10111011",	-- 0x026d
		"11001101",	-- 0x026e
		"10101010",	-- 0x026f
		"11100110",	-- 0x0270
		"10001111",	-- 0x0271
		"00001000",	-- 0x0272
		"00001010",	-- 0x0273
		"11111111",	-- 0x0274
		"00100000",	-- 0x0275
		"11001011",	-- 0x0276
		"00111100",	-- 0x0277
		"10100001",	-- 0x0278
		"01011010",	-- 0x0279
		"10100001",	-- 0x027a
		"10100000",	-- 0x027b
		"01111110",	-- 0x027c
		"00000100",	-- 0x027d
		"00101000",	-- 0x027e
		"11111010",	-- 0x027f
		"01010000",	-- 0x0280
		"01111101",	-- 0x0281
		"10100000",	-- 0x0282
		"01011110",	-- 0x0283
		"00001110",	-- 0x0284
		"00011111",	-- 0x0285
		"10101011",	-- 0x0286
		"00111110",	-- 0x0287
		"10011110",	-- 0x0288
		"01011101",	-- 0x0289
		"10010101",	-- 0x028a
		"01111100",	-- 0x028b
		"10000000",	-- 0x028c
		"10011100",	-- 0x028d
		"10000000",	-- 0x028e
		"10111100",	-- 0x028f
		"10000000",	-- 0x0290
		"11010010",	-- 0x0291
		"10000000",	-- 0x0292
		"11100100",	-- 0x0293
		"10000000",	-- 0x0294
		"00001110",	-- 0x0295
		"00011111",	-- 0x0296
		"10101011",	-- 0x0297
		"00111110",	-- 0x0298
		"10011110",	-- 0x0299
		"01011101",	-- 0x029a
		"10010101",	-- 0x029b
		"01111100",	-- 0x029c
		"10000000",	-- 0x029d
		"10011100",	-- 0x029e
		"01101011",	-- 0x029f
		"10111100",	-- 0x02a0
		"01101111",	-- 0x02a1
		"11010010",	-- 0x02a2
		"10000000",	-- 0x02a3
		"11100100",	-- 0x02a4
		"10000000",	-- 0x02a5
		"00001110",	-- 0x02a6
		"00011111",	-- 0x02a7
		"10101011",	-- 0x02a8
		"00111110",	-- 0x02a9
		"10011110",	-- 0x02aa
		"01011101",	-- 0x02ab
		"10010101",	-- 0x02ac
		"01111100",	-- 0x02ad
		"10000000",	-- 0x02ae
		"10011100",	-- 0x02af
		"10000000",	-- 0x02b0
		"10111100",	-- 0x02b1
		"10000000",	-- 0x02b2
		"11010010",	-- 0x02b3
		"10000000",	-- 0x02b4
		"11100100",	-- 0x02b5
		"10000000",	-- 0x02b6
		"00000000",	-- 0x02b7
		"11000000",	-- 0x02b8
		"00110011",	-- 0x02b9
		"01000000",	-- 0x02ba
		"01001000",	-- 0x02bb
		"01010101",	-- 0x02bc
		"01110011",	-- 0x02bd
		"01111011",	-- 0x02be
		"10001000",	-- 0x02bf
		"00001000",	-- 0x02c0
		"01100000",	-- 0x02c1
		"00000101",	-- 0x02c2
		"01010110",	-- 0x02c3
		"01010110",	-- 0x02c4
		"01101011",	-- 0x02c5
		"10000000",	-- 0x02c6
		"10010110",	-- 0x02c7
		"11001101",	-- 0x02c8
		"00000101",	-- 0x02c9
		"00010001",	-- 0x02ca
		"00000101",	-- 0x02cb
		"00010001",	-- 0x02cc
		"00011010",	-- 0x02cd
		"10000000",	-- 0x02ce
		"11001000",	-- 0x02cf
		"11001000",	-- 0x02d0
		"11001000",	-- 0x02d1
		"11001000",	-- 0x02d2
		"11001000",	-- 0x02d3
		"01010110",	-- 0x02d4
		"10000000",	-- 0x02d5
		"00000000",	-- 0x02d6
		"00001100",	-- 0x02d7
		"00101010",	-- 0x02d8
		"01000000",	-- 0x02d9
		"10010101",	-- 0x02da
		"00000000",	-- 0x02db
		"10000000",	-- 0x02dc
		"00000000",	-- 0x02dd
		"00011110",	-- 0x02de
		"00110011",	-- 0x02df
		"01000000",	-- 0x02e0
		"01000000",	-- 0x02e1
		"00000010",	-- 0x02e2
		"11010010",	-- 0x02e3
		"01000000",	-- 0x02e4
		"11100100",	-- 0x02e5
		"00000000",	-- 0x02e6
		"00011010",	-- 0x02e7
		"10000000",	-- 0x02e8
		"00000110",	-- 0x02e9
		"00001010",	-- 0x02ea
		"00011001",	-- 0x02eb
		"00100101",	-- 0x02ec
		"00100101",	-- 0x02ed
		"01001111",	-- 0x02ee
		"01000000",	-- 0x02ef
		"10000000",	-- 0x02f0
		"00000000",	-- 0x02f1
		"00100000",	-- 0x02f2
		"01000000",	-- 0x02f3
		"00101001",	-- 0x02f4
		"00111010",	-- 0x02f5
		"01001101",	-- 0x02f6
		"00000100",	-- 0x02f7
		"00101000",	-- 0x02f8
		"01000100",	-- 0x02f9
		"01010000",	-- 0x02fa
		"01000100",	-- 0x02fb
		"01111000",	-- 0x02fc
		"01000100",	-- 0x02fd
		"00000110",	-- 0x02fe
		"00000000",	-- 0x02ff
		"00000100",	-- 0x0300
		"00000010",	-- 0x0301
		"00000000",	-- 0x0302
		"00000100",	-- 0x0303
		"11010000",	-- 0x0304
		"11010000",	-- 0x0305
		"11010000",	-- 0x0306
		"11010000",	-- 0x0307
		"11010000",	-- 0x0308
		"10110110",	-- 0x0309
		"01101010",	-- 0x030a
		"01100100",	-- 0x030b
		"01011111",	-- 0x030c
		"01111001",	-- 0x030d
		"01011010",	-- 0x030e
		"01011010",	-- 0x030f
		"01010000",	-- 0x0310
		"01000110",	-- 0x0311
		"01000110",	-- 0x0312
		"01010000",	-- 0x0313
		"01010000",	-- 0x0314
		"01010000",	-- 0x0315
		"01000110",	-- 0x0316
		"00110001",	-- 0x0317
		"01000110",	-- 0x0318
		"00110001",	-- 0x0319
		"00110001",	-- 0x031a
		"00110001",	-- 0x031b
		"00110001",	-- 0x031c
		"01010000",	-- 0x031d
		"00110000",	-- 0x031e
		"00000000",	-- 0x031f
		"01100110",	-- 0x0320
		"10011010",	-- 0x0321
		"11001101",	-- 0x0322
		"00010010",	-- 0x0323
		"00100110",	-- 0x0324
		"01111010",	-- 0x0325
		"00111010",	-- 0x0326
		"01011111",	-- 0x0327
		"01010001",	-- 0x0328
		"01001111",	-- 0x0329
		"01101011",	-- 0x032a
		"01001000",	-- 0x032b
		"10000110",	-- 0x032c
		"00111101",	-- 0x032d
		"10110011",	-- 0x032e
		"00110011",	-- 0x032f
		"11010010",	-- 0x0330
		"00101001",	-- 0x0331
		"11011100",	-- 0x0332
		"00010110",	-- 0x0333
		"11100001",	-- 0x0334
		"00010001",	-- 0x0335
		"11100100",	-- 0x0336
		"00000000",	-- 0x0337
		"00001010",	-- 0x0338
		"00100110",	-- 0x0339
		"00010100",	-- 0x033a
		"00111010",	-- 0x033b
		"00010100",	-- 0x033c
		"01010001",	-- 0x033d
		"00010100",	-- 0x033e
		"10000110",	-- 0x033f
		"00010100",	-- 0x0340
		"11011100",	-- 0x0341
		"00010100",	-- 0x0342
		"11101000",	-- 0x0343
		"00011010",	-- 0x0344
		"00000010",	-- 0x0345
		"10110011",	-- 0x0346
		"00001010",	-- 0x0347
		"11010010",	-- 0x0348
		"00110011",	-- 0x0349
		"00011111",	-- 0x034a
		"00001010",	-- 0x034b
		"00100001",	-- 0x034c
		"00110000",	-- 0x034d
		"00000000",	-- 0x034e
		"00100110",	-- 0x034f
		"00100110",	-- 0x0350
		"00100110",	-- 0x0351
		"00011010",	-- 0x0352
		"00100000",	-- 0x0353
		"10010010",	-- 0x0354
		"01000000",	-- 0x0355
		"00000000",	-- 0x0356
		"00000000",	-- 0x0357
		"01101010",	-- 0x0358
		"01111010",	-- 0x0359
		"10000101",	-- 0x035a
		"10010101",	-- 0x035b
		"11111111",	-- 0x035c
		"10000011",	-- 0x035d
		"10000001",	-- 0x035e
		"10000000",	-- 0x035f
		"01111111",	-- 0x0360
		"01111101",	-- 0x0361
		"01101010",	-- 0x0362
		"01111010",	-- 0x0363
		"10000101",	-- 0x0364
		"10010101",	-- 0x0365
		"11111111",	-- 0x0366
		"10000011",	-- 0x0367
		"10000001",	-- 0x0368
		"10000000",	-- 0x0369
		"01111111",	-- 0x036a
		"01111101",	-- 0x036b
		"01110000",	-- 0x036c
		"10010000",	-- 0x036d
		"10100000",	-- 0x036e
		"10110000",	-- 0x036f
		"01110000",	-- 0x0370
		"10010000",	-- 0x0371
		"00010000",	-- 0x0372
		"00000000",	-- 0x0373
		"00000000",	-- 0x0374
		"00000000",	-- 0x0375
		"00001100",	-- 0x0376
		"00100110",	-- 0x0377
		"11110011",	-- 0x0378
		"01010001",	-- 0x0379
		"11110001",	-- 0x037a
		"01101011",	-- 0x037b
		"11101000",	-- 0x037c
		"10000110",	-- 0x037d
		"11010111",	-- 0x037e
		"10110011",	-- 0x037f
		"10101100",	-- 0x0380
		"11010010",	-- 0x0381
		"10010100",	-- 0x0382
		"11100100",	-- 0x0383
		"10001101",	-- 0x0384
		"01110011",	-- 0x0385
		"01100000",	-- 0x0386
		"00011001",	-- 0x0387
		"00100111",	-- 0x0388
		"00110011",	-- 0x0389
		"00111011",	-- 0x038a
		"01110011",	-- 0x038b
		"01100000",	-- 0x038c
		"00110110",	-- 0x038d
		"00110011",	-- 0x038e
		"00110001",	-- 0x038f
		"00101100",	-- 0x0390
		"00000000",	-- 0x0391
		"00001000",	-- 0x0392
		"00010000",	-- 0x0393
		"00100000",	-- 0x0394
		"00000010",	-- 0x0395
		"00000100",	-- 0x0396
		"00000110",	-- 0x0397
		"00000001",	-- 0x0398
		"00000001",	-- 0x0399
		"00000010",	-- 0x039a
		"01110000",	-- 0x039b
		"11000000",	-- 0x039c
		"01101000",	-- 0x039d
		"11000000",	-- 0x039e
		"01101000",	-- 0x039f
		"10111000",	-- 0x03a0
		"11100110",	-- 0x03a1
		"00000000",	-- 0x03a2
		"00011010",	-- 0x03a3
		"00000000",	-- 0x03a4
		"11100110",	-- 0x03a5
		"00011010",	-- 0x03a6
		"11100110",	-- 0x03a7
		"00011010",	-- 0x03a8
		"11100110",	-- 0x03a9
		"00011010",	-- 0x03aa
		"11100110",	-- 0x03ab
		"00011010",	-- 0x03ac
		"11100110",	-- 0x03ad
		"00011010",	-- 0x03ae
		"11100110",	-- 0x03af
		"00011010",	-- 0x03b0
		"11100110",	-- 0x03b1
		"00011010",	-- 0x03b2
		"11100110",	-- 0x03b3
		"00011010",	-- 0x03b4
		"10101110",	-- 0x03b5
		"01010010",	-- 0x03b6
		"10000000",	-- 0x03b7
		"00000000",	-- 0x03b8
		"01110101",	-- 0x03b9
		"00110000",	-- 0x03ba
		"00000000",	-- 0x03bb
		"10101111",	-- 0x03bc
		"01100100",	-- 0x03bd
		"00110111",	-- 0x03be
		"10001000",	-- 0x03bf
		"00101010",	-- 0x03c0
		"00000101",	-- 0x03c1
		"00000000",	-- 0x03c2
		"00000000",	-- 0x03c3
		"00000000",	-- 0x03c4
		"01111000",	-- 0x03c5
		"01000101",	-- 0x03c6
		"11100110",	-- 0x03c7
		"00011010",	-- 0x03c8
		"11111100",	-- 0x03c9
		"00000111",	-- 0x03ca
		"11111100",	-- 0x03cb
		"00000111",	-- 0x03cc
		"11111100",	-- 0x03cd
		"00000111",	-- 0x03ce
		"11111011",	-- 0x03cf
		"00001101",	-- 0x03d0
		"00110001",	-- 0x03d1
		"00000101",	-- 0x03d2
		"11000011",	-- 0x03d3
		"00010100",	-- 0x03d4
		"11000011",	-- 0x03d5
		"00010100",	-- 0x03d6
		"00011111",	-- 0x03d7
		"11101101",	-- 0x03d8
		"10000001",	-- 0x03d9
		"01000010",	-- 0x03da
		"00001110",	-- 0x03db
		"11101010",	-- 0x03dc
		"10000001",	-- 0x03dd
		"01000000",	-- 0x03de
		"00000101",	-- 0x03df
		"10101001",	-- 0x03e0
		"10000000",	-- 0x03e1
		"01000010",	-- 0x03e2
		"00000110",	-- 0x03e3
		"00011101",	-- 0x03e4
		"00011101",	-- 0x03e5
		"10101001",	-- 0x03e6
		"10000000",	-- 0x03e7
		"01000100",	-- 0x03e8
		"00000011",	-- 0x03e9
		"10100110",	-- 0x03ea
		"10000000",	-- 0x03eb
		"01100111",	-- 0x03ec
		"01100011",	-- 0x03ed
		"11011010",	-- 0x03ee
		"01010111",	-- 0x03ef
		"01010011",	-- 0x03f0
		"10001100",	-- 0x03f1
		"10010110",	-- 0x03f2
		"01011001",	-- 0x03f3
		"00111110",	-- 0x03f4
		"00011010",	-- 0x03f5
		"01101111",	-- 0x03f6
		"00001101",	-- 0x03f7
		"00111100",	-- 0x03f8
		"11101100",	-- 0x03f9
		"10000000",	-- 0x03fa
		"01000101",	-- 0x03fb
		"00000011",	-- 0x03fc
		"01111110",	-- 0x03fd
		"01000000",	-- 0x03fe
		"00000101",	-- 0x03ff
		"01111111",	-- 0x0400
		"11101100",	-- 0x0401
		"10000000",	-- 0x0402
		"01000100",	-- 0x0403
		"00000110",	-- 0x0404
		"11101010",	-- 0x0405
		"10000001",	-- 0x0406
		"01010011",	-- 0x0407
		"01100011",	-- 0x0408
		"00011101",	-- 0x0409
		"00011101",	-- 0x040a
		"11101100",	-- 0x040b
		"10000010",	-- 0x040c
		"01000100",	-- 0x040d
		"11111010",	-- 0x040e
		"11101010",	-- 0x040f
		"10000010",	-- 0x0410
		"11100100",	-- 0x0411
		"10000000",	-- 0x0412
		"01101100",	-- 0x0413
		"00111100",	-- 0x0414
		"11100100",	-- 0x0415
		"10000000",	-- 0x0416
		"00101110",	-- 0x0417
		"10100101",	-- 0x0418
		"00000000",	-- 0x0419
		"00101101",	-- 0x041a
		"11101010",	-- 0x041b
		"10000011",	-- 0x041c
		"11100100",	-- 0x041d
		"10000001",	-- 0x041e
		"01000100",	-- 0x041f
		"00000110",	-- 0x0420
		"01010100",	-- 0x0421
		"01010101",	-- 0x0422
		"01000111",	-- 0x0423
		"11100000",	-- 0x0424
		"00011101",	-- 0x0425
		"00011101",	-- 0x0426
		"01101101",	-- 0x0427
		"00101110",	-- 0x0428
		"10100001",	-- 0x0429
		"00000000",	-- 0x042a
		"11100000",	-- 0x042b
		"10000001",	-- 0x042c
		"00101101",	-- 0x042d
		"01100011",	-- 0x042e
		"00000100",	-- 0x042f
		"00000100",	-- 0x0430
		"00000100",	-- 0x0431
		"00000100",	-- 0x0432
		"00000100",	-- 0x0433
		"01000000",	-- 0x0434
		"00000010",	-- 0x0435
		"00000110",	-- 0x0436
		"00000110",	-- 0x0437
		"01100001",	-- 0x0438
		"00111100",	-- 0x0439
		"01000000",	-- 0x043a
		"00011101",	-- 0x043b
		"11011011",	-- 0x043c
		"01010111",	-- 0x043d
		"11001010",	-- 0x043e
		"00000100",	-- 0x043f
		"01000000",	-- 0x0440
		"00000111",	-- 0x0441
		"11011011",	-- 0x0442
		"01010111",	-- 0x0443
		"11001010",	-- 0x0444
		"00001000",	-- 0x0445
		"10001100",	-- 0x0446
		"11001010",	-- 0x0447
		"00010000",	-- 0x0448
		"11100101",	-- 0x0449
		"10000000",	-- 0x044a
		"01000101",	-- 0x044b
		"00100101",	-- 0x044c
		"01101100",	-- 0x044d
		"11101101",	-- 0x044e
		"10000001",	-- 0x044f
		"01000011",	-- 0x0450
		"00000010",	-- 0x0451
		"11101011",	-- 0x0452
		"10000001",	-- 0x0453
		"00101110",	-- 0x0454
		"01011010",	-- 0x0455
		"10100001",	-- 0x0456
		"00000000",	-- 0x0457
		"00101101",	-- 0x0458
		"11000000",	-- 0x0459
		"00000010",	-- 0x045a
		"00001101",	-- 0x045b
		"01011010",	-- 0x045c
		"01000111",	-- 0x045d
		"00010000",	-- 0x045e
		"01101101",	-- 0x045f
		"00101110",	-- 0x0460
		"11101010",	-- 0x0461
		"10000001",	-- 0x0462
		"11100100",	-- 0x0463
		"10000000",	-- 0x0464
		"01000100",	-- 0x0465
		"00000101",	-- 0x0466
		"01010100",	-- 0x0467
		"01010101",	-- 0x0468
		"01101011",	-- 0x0469
		"00000000",	-- 0x046a
		"00011101",	-- 0x046b
		"10100001",	-- 0x046c
		"00000000",	-- 0x046d
		"00101101",	-- 0x046e
		"11100000",	-- 0x046f
		"10000000",	-- 0x0470
		"01100011",	-- 0x0471
		"11101010",	-- 0x0472
		"10000010",	-- 0x0473
		"01010011",	-- 0x0474
		"01100011",	-- 0x0475
		"10101000",	-- 0x0476
		"10000000",	-- 0x0477
		"01000100",	-- 0x0478
		"00000010",	-- 0x0479
		"01010010",	-- 0x047a
		"01010011",	-- 0x047b
		"11101100",	-- 0x047c
		"10000010",	-- 0x047d
		"01000101",	-- 0x047e
		"00000011",	-- 0x047f
		"11101010",	-- 0x0480
		"10000010",	-- 0x0481
		"01010011",	-- 0x0482
		"00011101",	-- 0x0483
		"01100011",	-- 0x0484
		"00000100",	-- 0x0485
		"00000100",	-- 0x0486
		"00000100",	-- 0x0487
		"00000100",	-- 0x0488
		"00000100",	-- 0x0489
		"01100001",	-- 0x048a
		"11101010",	-- 0x048b
		"01101110",	-- 0x048c
		"10011010",	-- 0x048d
		"01111000",	-- 0x048e
		"00111101",	-- 0x048f
		"00111110",	-- 0x0490
		"00011101",	-- 0x0491
		"00011101",	-- 0x0492
		"01111000",	-- 0x0493
		"01100001",	-- 0x0494
		"11100000",	-- 0x0495
		"01101101",	-- 0x0496
		"11101011",	-- 0x0497
		"00000001",	-- 0x0498
		"01010111",	-- 0x0499
		"01101101",	-- 0x049a
		"00101110",	-- 0x049b
		"10100001",	-- 0x049c
		"00000000",	-- 0x049d
		"00111011",	-- 0x049e
		"01111010",	-- 0x049f
		"10010111",	-- 0x04a0
		"01111010",	-- 0x04a1
		"00111111",	-- 0x04a2
		"01101111",	-- 0x04a3
		"10010110",	-- 0x04a4
		"01111000",	-- 0x04a5
		"01100001",	-- 0x04a6
		"10110001",	-- 0x04a7
		"10010010",	-- 0x04a8
		"01111010",	-- 0x04a9
		"01111111",	-- 0x04aa
		"01111101",	-- 0x04ab
		"00001111",	-- 0x04ac
		"10010110",	-- 0x04ad
		"01111000",	-- 0x04ae
		"01100001",	-- 0x04af
		"10101000",	-- 0x04b0
		"10010010",	-- 0x04b1
		"01111011",	-- 0x04b2
		"10001111",	-- 0x04b3
		"00000000",	-- 0x04b4
		"01111010",	-- 0x04b5
		"01111101",	-- 0x04b6
		"01000000",	-- 0x04b7
		"10100011",	-- 0x04b8
		"10001110",	-- 0x04b9
		"00000000",	-- 0x04ba
		"00000000",	-- 0x04bb
		"00001100",	-- 0x04bc
		"11101010",	-- 0x04bd
		"00000000",	-- 0x04be
		"01010110",	-- 0x04bf
		"01000111",	-- 0x04c0
		"00000010",	-- 0x04c1
		"01100110",	-- 0x04c2
		"00000000",	-- 0x04c3
		"00011100",	-- 0x04c4
		"01010001",	-- 0x04c5
		"01000110",	-- 0x04c6
		"11110101",	-- 0x04c7
		"01100011",	-- 0x04c8
		"00000100",	-- 0x04c9
		"00000100",	-- 0x04ca
		"00000100",	-- 0x04cb
		"00000100",	-- 0x04cc
		"00000100",	-- 0x04cd
		"00000100",	-- 0x04ce
		"00000100",	-- 0x04cf
		"01100011",	-- 0x04d0
		"00011000",	-- 0x04d1
		"00010101",	-- 0x04d2
		"00011000",	-- 0x04d3
		"00010101",	-- 0x04d4
		"00011000",	-- 0x04d5
		"00010101",	-- 0x04d6
		"00011000",	-- 0x04d7
		"00010101",	-- 0x04d8
		"01100011",	-- 0x04d9
		"00000100",	-- 0x04da
		"00000100",	-- 0x04db
		"00000100",	-- 0x04dc
		"00000100",	-- 0x04dd
		"00000100",	-- 0x04de
		"00000100",	-- 0x04df
		"00000100",	-- 0x04e0
		"01011000",	-- 0x04e1
		"01000111",	-- 0x04e2
		"00000010",	-- 0x04e3
		"11001011",	-- 0x04e4
		"11111111",	-- 0x04e5
		"01100011",	-- 0x04e6
		"01110111",	-- 0x04e7
		"00011000",	-- 0x04e8
		"00110111",	-- 0x04e9
		"00011000",	-- 0x04ea
		"00000100",	-- 0x04eb
		"01010100",	-- 0x04ec
		"01010101",	-- 0x04ed
		"10000100",	-- 0x04ee
		"00000000",	-- 0x04ef
		"01100011",	-- 0x04f0
		"01010010",	-- 0x04f1
		"10000111",	-- 0x04f2
		"00000001",	-- 0x04f3
		"10000000",	-- 0x04f4
		"01100001",	-- 0x04f5
		"00010000",	-- 0x04f6
		"00111101",	-- 0x04f7
		"01101100",	-- 0x04f8
		"00111100",	-- 0x04f9
		"00000100",	-- 0x04fa
		"11000010",	-- 0x04fb
		"11111111",	-- 0x04fc
		"01111100",	-- 0x04fd
		"01000111",	-- 0x04fe
		"00000100",	-- 0x04ff
		"10000110",	-- 0x0500
		"11111111",	-- 0x0501
		"11111111",	-- 0x0502
		"01100111",	-- 0x0503
		"00000010",	-- 0x0504
		"00010101",	-- 0x0505
		"01100011",	-- 0x0506
		"01101000",	-- 0x0507
		"01101110",	-- 0x0508
		"00101110",	-- 0x0509
		"10100001",	-- 0x050a
		"00000000",	-- 0x050b
		"00111111",	-- 0x050c
		"11101010",	-- 0x050d
		"00000000",	-- 0x050e
		"10100001",	-- 0x050f
		"00000011",	-- 0x0510
		"00001101",	-- 0x0511
		"10100011",	-- 0x0512
		"00000000",	-- 0x0513
		"11101010",	-- 0x0514
		"00000001",	-- 0x0515
		"10100001",	-- 0x0516
		"00000011",	-- 0x0517
		"10100011",	-- 0x0518
		"00000011",	-- 0x0519
		"01101010",	-- 0x051a
		"00000010",	-- 0x051b
		"10100001",	-- 0x051c
		"00000001",	-- 0x051d
		"11100001",	-- 0x051e
		"00000000",	-- 0x051f
		"10000000",	-- 0x0520
		"00000000",	-- 0x0521
		"00001101",	-- 0x0522
		"01010010",	-- 0x0523
		"11100001",	-- 0x0524
		"00000010",	-- 0x0525
		"00010110",	-- 0x0526
		"00001101",	-- 0x0527
		"10100011",	-- 0x0528
		"00000010",	-- 0x0529
		"00101011",	-- 0x052a
		"00000000",	-- 0x052b
		"11101010",	-- 0x052c
		"00000000",	-- 0x052d
		"01000111",	-- 0x052e
		"00000100",	-- 0x052f
		"10000110",	-- 0x0530
		"11111111",	-- 0x0531
		"11111111",	-- 0x0532
		"10001100",	-- 0x0533
		"10100110",	-- 0x0534
		"00000001",	-- 0x0535
		"01111110",	-- 0x0536
		"01111111",	-- 0x0537
		"01100011",	-- 0x0538
		"00111100",	-- 0x0539
		"11001110",	-- 0x053a
		"11111000",	-- 0x053b
		"01000111",	-- 0x053c
		"00000100",	-- 0x053d
		"10000110",	-- 0x053e
		"01111111",	-- 0x053f
		"11111111",	-- 0x0540
		"01100011",	-- 0x0541
		"00000110",	-- 0x0542
		"00000110",	-- 0x0543
		"00000110",	-- 0x0544
		"00000110",	-- 0x0545
		"00000110",	-- 0x0546
		"00111110",	-- 0x0547
		"00111101",	-- 0x0548
		"10000001",	-- 0x0549
		"00100000",	-- 0x054a
		"00001100",	-- 0x054b
		"00111100",	-- 0x054c
		"00000100",	-- 0x054d
		"01100011",	-- 0x054e
		"01100001",	-- 0x054f
		"00001001",	-- 0x0550
		"00010111",	-- 0x0551
		"00010110",	-- 0x0552
		"01000100",	-- 0x0553
		"00000011",	-- 0x0554
		"10000110",	-- 0x0555
		"11111111",	-- 0x0556
		"11111111",	-- 0x0557
		"00111110",	-- 0x0558
		"01100011",	-- 0x0559
		"01011010",	-- 0x055a
		"01101110",	-- 0x055b
		"00101110",	-- 0x055c
		"01101010",	-- 0x055d
		"00000001",	-- 0x055e
		"10100001",	-- 0x055f
		"00000001",	-- 0x0560
		"01101101",	-- 0x0561
		"01101010",	-- 0x0562
		"00000001",	-- 0x0563
		"10100001",	-- 0x0564
		"00000000",	-- 0x0565
		"00111110",	-- 0x0566
		"01111000",	-- 0x0567
		"01111101",	-- 0x0568
		"00001110",	-- 0x0569
		"00010010",	-- 0x056a
		"00111100",	-- 0x056b
		"01100011",	-- 0x056c
		"01101101",	-- 0x056d
		"00111100",	-- 0x056e
		"10101000",	-- 0x056f
		"10000000",	-- 0x0570
		"01000111",	-- 0x0571
		"00100101",	-- 0x0572
		"01000100",	-- 0x0573
		"00010100",	-- 0x0574
		"01010100",	-- 0x0575
		"01010101",	-- 0x0576
		"10000100",	-- 0x0577
		"00000000",	-- 0x0578
		"00111110",	-- 0x0579
		"01111100",	-- 0x057a
		"01100001",	-- 0x057b
		"11011110",	-- 0x057c
		"10001001",	-- 0x057d
		"00000000",	-- 0x057e
		"00000000",	-- 0x057f
		"01000110",	-- 0x0580
		"00000001",	-- 0x0581
		"01010111",	-- 0x0582
		"01010100",	-- 0x0583
		"01010101",	-- 0x0584
		"10000100",	-- 0x0585
		"00000000",	-- 0x0586
		"01000000",	-- 0x0587
		"00001010",	-- 0x0588
		"00111110",	-- 0x0589
		"01111100",	-- 0x058a
		"01100001",	-- 0x058b
		"11001110",	-- 0x058c
		"10001001",	-- 0x058d
		"00000000",	-- 0x058e
		"00000000",	-- 0x058f
		"01000110",	-- 0x0590
		"00000001",	-- 0x0591
		"01010111",	-- 0x0592
		"10100111",	-- 0x0593
		"10000000",	-- 0x0594
		"10101010",	-- 0x0595
		"10000000",	-- 0x0596
		"10001100",	-- 0x0597
		"00101101",	-- 0x0598
		"00111100",	-- 0x0599
		"01100011",	-- 0x059a
		"10001111",	-- 0x059b
		"11111111",	-- 0x059c
		"11111000",	-- 0x059d
		"01101000",	-- 0x059e
		"00111100",	-- 0x059f
		"10001001",	-- 0x05a0
		"00000000",	-- 0x05a1
		"00000000",	-- 0x05a2
		"01000110",	-- 0x05a3
		"00000101",	-- 0x05a4
		"01111110",	-- 0x05a5
		"01000000",	-- 0x05a6
		"01011001",	-- 0x05a7
		"00011111",	-- 0x05a8
		"00000110",	-- 0x05a9
		"01001010",	-- 0x05aa
		"11111100",	-- 0x05ab
		"00011101",	-- 0x05ac
		"00000100",	-- 0x05ad
		"00111110",	-- 0x05ae
		"01111000",	-- 0x05af
		"10001001",	-- 0x05b0
		"00000000",	-- 0x05b1
		"00000000",	-- 0x05b2
		"01000111",	-- 0x05b3
		"01000111",	-- 0x05b4
		"01001011",	-- 0x05b5
		"00000100",	-- 0x05b6
		"00011101",	-- 0x05b7
		"00000110",	-- 0x05b8
		"01001010",	-- 0x05b9
		"11111100",	-- 0x05ba
		"01101111",	-- 0x05bb
		"01101001",	-- 0x05bc
		"01010110",	-- 0x05bd
		"01101000",	-- 0x05be
		"01101111",	-- 0x05bf
		"00101110",	-- 0x05c0
		"01000111",	-- 0x05c1
		"00001010",	-- 0x05c2
		"00111101",	-- 0x05c3
		"10100101",	-- 0x05c4
		"00000010",	-- 0x05c5
		"10100011",	-- 0x05c6
		"00000000",	-- 0x05c7
		"01010011",	-- 0x05c8
		"10100101",	-- 0x05c9
		"00000010",	-- 0x05ca
		"10100011",	-- 0x05cb
		"00000001",	-- 0x05cc
		"00111101",	-- 0x05cd
		"01100000",	-- 0x05ce
		"00000010",	-- 0x05cf
		"10100101",	-- 0x05d0
		"00000010",	-- 0x05d1
		"01101101",	-- 0x05d2
		"01010011",	-- 0x05d3
		"10100101",	-- 0x05d4
		"00000010",	-- 0x05d5
		"01111100",	-- 0x05d6
		"01100100",	-- 0x05d7
		"00000011",	-- 0x05d8
		"01000111",	-- 0x05d9
		"00001101",	-- 0x05da
		"10101000",	-- 0x05db
		"00000000",	-- 0x05dc
		"01101101",	-- 0x05dd
		"10100001",	-- 0x05de
		"00000011",	-- 0x05df
		"00111111",	-- 0x05e0
		"01111100",	-- 0x05e1
		"10100001",	-- 0x05e2
		"00000011",	-- 0x05e3
		"00001101",	-- 0x05e4
		"00111101",	-- 0x05e5
		"10100111",	-- 0x05e6
		"00000000",	-- 0x05e7
		"01111110",	-- 0x05e8
		"01111110",	-- 0x05e9
		"01111111",	-- 0x05ea
		"10001101",	-- 0x05eb
		"00000000",	-- 0x05ec
		"00000000",	-- 0x05ed
		"01001010",	-- 0x05ee
		"00000100",	-- 0x05ef
		"00000100",	-- 0x05f0
		"00011101",	-- 0x05f1
		"01001011",	-- 0x05f2
		"11111100",	-- 0x05f3
		"01000111",	-- 0x05f4
		"00001011",	-- 0x05f5
		"00000110",	-- 0x05f6
		"01000101",	-- 0x05f7
		"00000011",	-- 0x05f8
		"00011111",	-- 0x05f9
		"01000000",	-- 0x05fa
		"11111000",	-- 0x05fb
		"10000110",	-- 0x05fc
		"11111111",	-- 0x05fd
		"11111111",	-- 0x05fe
		"01100111",	-- 0x05ff
		"01000001",	-- 0x0600
		"01100101",	-- 0x0601
		"01100011",	-- 0x0602
		"00110011",	-- 0x0603
		"00000111",	-- 0x0604
		"00011111",	-- 0x0605
		"00000101",	-- 0x0606
		"00110011",	-- 0x0607
		"00011000",	-- 0x0608
		"00010000",	-- 0x0609
		"00110011",	-- 0x060a
		"00000000",	-- 0x060b
		"00011101",	-- 0x060c
		"00110011",	-- 0x060d
		"00110000",	-- 0x060e
		"00010011",	-- 0x060f
		"00110011",	-- 0x0610
		"11110100",	-- 0x0611
		"00010010",	-- 0x0612
		"00110011",	-- 0x0613
		"11111001",	-- 0x0614
		"00000011",	-- 0x0615
		"10000110",	-- 0x0616
		"10000001",	-- 0x0617
		"11011110",	-- 0x0618
		"10011010",	-- 0x0619
		"00011000",	-- 0x061a
		"10000110",	-- 0x061b
		"10010010",	-- 0x061c
		"00000000",	-- 0x061d
		"10011010",	-- 0x061e
		"00011010",	-- 0x061f
		"00110011",	-- 0x0620
		"11111100",	-- 0x0621
		"00010100",	-- 0x0622
		"00110011",	-- 0x0623
		"00110000",	-- 0x0624
		"00000111",	-- 0x0625
		"00110011",	-- 0x0626
		"11011101",	-- 0x0627
		"00100000",	-- 0x0628
		"01110010",	-- 0x0629
		"00100001",	-- 0x062a
		"00110011",	-- 0x062b
		"11011001",	-- 0x062c
		"00100010",	-- 0x062d
		"01110010",	-- 0x062e
		"00100011",	-- 0x062f
		"00110011",	-- 0x0630
		"00000011",	-- 0x0631
		"00101001",	-- 0x0632
		"10000110",	-- 0x0633
		"00000001",	-- 0x0634
		"00000111",	-- 0x0635
		"10011010",	-- 0x0636
		"00000000",	-- 0x0637
		"00110011",	-- 0x0638
		"11100011",	-- 0x0639
		"00010001",	-- 0x063a
		"00110011",	-- 0x063b
		"00111111",	-- 0x063c
		"00100100",	-- 0x063d
		"11011010",	-- 0x063e
		"00101001",	-- 0x063f
		"11000010",	-- 0x0640
		"10000000",	-- 0x0641
		"00010000",	-- 0x0642
		"00010000",	-- 0x0643
		"11011000",	-- 0x0644
		"00100100",	-- 0x0645
		"10010010",	-- 0x0646
		"00100100",	-- 0x0647
		"00110011",	-- 0x0648
		"00000000",	-- 0x0649
		"00100110",	-- 0x064a
		"00110011",	-- 0x064b
		"00000000",	-- 0x064c
		"00100111",	-- 0x064d
		"01110111",	-- 0x064e
		"01001011",	-- 0x064f
		"11011010",	-- 0x0650
		"00101011",	-- 0x0651
		"11011010",	-- 0x0652
		"00000110",	-- 0x0653
		"01110101",	-- 0x0654
		"01101011",	-- 0x0655
		"01110111",	-- 0x0656
		"00101011",	-- 0x0657
		"00110011",	-- 0x0658
		"10010000",	-- 0x0659
		"00000110",	-- 0x065a
		"01010010",	-- 0x065b
		"01010011",	-- 0x065c
		"10011010",	-- 0x065d
		"00101100",	-- 0x065e
		"10011010",	-- 0x065f
		"00101110",	-- 0x0660
		"01110111",	-- 0x0661
		"01100110",	-- 0x0662
		"10001011",	-- 0x0663
		"00000010",	-- 0x0664
		"11111111",	-- 0x0665
		"01010010",	-- 0x0666
		"01010011",	-- 0x0667
		"10001111",	-- 0x0668
		"00000000",	-- 0x0669
		"01000000",	-- 0x066a
		"10000010",	-- 0x066b
		"10001101",	-- 0x066c
		"00000000",	-- 0x066d
		"01111111",	-- 0x066e
		"01000011",	-- 0x066f
		"11111010",	-- 0x0670
		"10001111",	-- 0x0671
		"00000000",	-- 0x0672
		"10100000",	-- 0x0673
		"10001010",	-- 0x0674
		"10001101",	-- 0x0675
		"00000010",	-- 0x0676
		"01000111",	-- 0x0677
		"01000011",	-- 0x0678
		"11111010",	-- 0x0679
		"00000001",	-- 0x067a
		"11110000",	-- 0x067b
		"00100000",	-- 0x067c
		"01110111",	-- 0x067d
		"00010110",	-- 0x067e
		"01110111",	-- 0x067f
		"10110000",	-- 0x0680
		"00110011",	-- 0x0681
		"11111111",	-- 0x0682
		"10110001",	-- 0x0683
		"00110011",	-- 0x0684
		"11111111",	-- 0x0685
		"11010111",	-- 0x0686
		"01110111",	-- 0x0687
		"01110010",	-- 0x0688
		"01110111",	-- 0x0689
		"01010010",	-- 0x068a
		"00110011",	-- 0x068b
		"11111111",	-- 0x068c
		"11000111",	-- 0x068d
		"01110111",	-- 0x068e
		"11010010",	-- 0x068f
		"00110011",	-- 0x0690
		"00000000",	-- 0x0691
		"01000001",	-- 0x0692
		"11001010",	-- 0x0693
		"00010000",	-- 0x0694
		"10110010",	-- 0x0695
		"00000001",	-- 0x0696
		"00000001",	-- 0x0697
		"00110011",	-- 0x0698
		"11111111",	-- 0x0699
		"10110011",	-- 0x069a
		"00110011",	-- 0x069b
		"11111111",	-- 0x069c
		"10110110",	-- 0x069d
		"00110011",	-- 0x069e
		"11111111",	-- 0x069f
		"10110111",	-- 0x06a0
		"11001010",	-- 0x06a1
		"01111000",	-- 0x06a2
		"10110010",	-- 0x06a3
		"00000001",	-- 0x06a4
		"01001000",	-- 0x06a5
		"10000110",	-- 0x06a6
		"00000000",	-- 0x06a7
		"10000000",	-- 0x06a8
		"10011010",	-- 0x06a9
		"01101011",	-- 0x06aa
		"00110011",	-- 0x06ab
		"10000000",	-- 0x06ac
		"01100000",	-- 0x06ad
		"00110011",	-- 0x06ae
		"11111111",	-- 0x06af
		"10101010",	-- 0x06b0
		"11001010",	-- 0x06b1
		"10000000",	-- 0x06b2
		"10110010",	-- 0x06b3
		"00000001",	-- 0x06b4
		"00011100",	-- 0x06b5
		"10000110",	-- 0x06b6
		"11001100",	-- 0x06b7
		"11001101",	-- 0x06b8
		"10111010",	-- 0x06b9
		"00000001",	-- 0x06ba
		"11000110",	-- 0x06bb
		"10000110",	-- 0x06bc
		"00000000",	-- 0x06bd
		"00000000",	-- 0x06be
		"10111010",	-- 0x06bf
		"00000001",	-- 0x06c0
		"11001000",	-- 0x06c1
		"00110011",	-- 0x06c2
		"11111110",	-- 0x06c3
		"11000100",	-- 0x06c4
		"00110011",	-- 0x06c5
		"11111110",	-- 0x06c6
		"11000101",	-- 0x06c7
		"11001010",	-- 0x06c8
		"11110100",	-- 0x06c9
		"10110010",	-- 0x06ca
		"00000001",	-- 0x06cb
		"11011101",	-- 0x06cc
		"01110111",	-- 0x06cd
		"01010101",	-- 0x06ce
		"11001010",	-- 0x06cf
		"11111110",	-- 0x06d0
		"10110010",	-- 0x06d1
		"00000001",	-- 0x06d2
		"01011010",	-- 0x06d3
		"11001010",	-- 0x06d4
		"11111111",	-- 0x06d5
		"10010010",	-- 0x06d6
		"10100110",	-- 0x06d7
		"11001010",	-- 0x06d8
		"11111111",	-- 0x06d9
		"10110010",	-- 0x06da
		"00000001",	-- 0x06db
		"01011101",	-- 0x06dc
		"10110010",	-- 0x06dd
		"00000001",	-- 0x06de
		"01011110",	-- 0x06df
		"10110010",	-- 0x06e0
		"00000001",	-- 0x06e1
		"01011111",	-- 0x06e2
		"11001010",	-- 0x06e3
		"10000000",	-- 0x06e4
		"10110010",	-- 0x06e5
		"00000001",	-- 0x06e6
		"01010110",	-- 0x06e7
		"01110000",	-- 0x06e8
		"10101001",	-- 0x06e9
		"11001010",	-- 0x06ea
		"11111111",	-- 0x06eb
		"10110010",	-- 0x06ec
		"00000001",	-- 0x06ed
		"10000111",	-- 0x06ee
		"11001010",	-- 0x06ef
		"11110011",	-- 0x06f0
		"10110010",	-- 0x06f1
		"00000001",	-- 0x06f2
		"10010100",	-- 0x06f3
		"10000110",	-- 0x06f4
		"00001000",	-- 0x06f5
		"10100100",	-- 0x06f6
		"10111010",	-- 0x06f7
		"00000001",	-- 0x06f8
		"10100001",	-- 0x06f9
		"10000110",	-- 0x06fa
		"00000100",	-- 0x06fb
		"00000000",	-- 0x06fc
		"10111010",	-- 0x06fd
		"00000001",	-- 0x06fe
		"10101111",	-- 0x06ff
		"11011010",	-- 0x0700
		"10011010",	-- 0x0701
		"10110010",	-- 0x0702
		"00000001",	-- 0x0703
		"10001110",	-- 0x0704
		"01010010",	-- 0x0705
		"01010011",	-- 0x0706
		"10011010",	-- 0x0707
		"00101100",	-- 0x0708
		"10000110",	-- 0x0709
		"00000000",	-- 0x070a
		"00001000",	-- 0x070b
		"10011010",	-- 0x070c
		"00101110",	-- 0x070d
		"00000111",	-- 0x070e
		"01010010",	-- 0x070f
		"10010010",	-- 0x0710
		"11111101",	-- 0x0711
		"01110111",	-- 0x0712
		"00101011",	-- 0x0713
		"01100111",	-- 0x0714
		"00010110",	-- 0x0715
		"10010010",	-- 0x0716
		"00000110",	-- 0x0717
		"00110111",	-- 0x0718
		"00110010",	-- 0x0719
		"11111101",	-- 0x071a
		"00000001",	-- 0x071b
		"11111011",	-- 0x071c
		"00011101",	-- 0x071d
		"00000001",	-- 0x071e
		"11111011",	-- 0x071f
		"00011101",	-- 0x0720
		"00000001",	-- 0x0721
		"11111001",	-- 0x0722
		"00100010",	-- 0x0723
		"01010010",	-- 0x0724
		"01010011",	-- 0x0725
		"10011010",	-- 0x0726
		"00101100",	-- 0x0727
		"10000110",	-- 0x0728
		"00000000",	-- 0x0729
		"00000100",	-- 0x072a
		"10011010",	-- 0x072b
		"00101110",	-- 0x072c
		"00000111",	-- 0x072d
		"00000001",	-- 0x072e
		"11111000",	-- 0x072f
		"01111100",	-- 0x0730
		"00000001",	-- 0x0731
		"11011111",	-- 0x0732
		"10100011",	-- 0x0733
		"00110101",	-- 0x0734
		"10111001",	-- 0x0735
		"00001011",	-- 0x0736
		"00110111",	-- 0x0737
		"11011001",	-- 0x0738
		"00001000",	-- 0x0739
		"01110111",	-- 0x073a
		"01010000",	-- 0x073b
		"11011010",	-- 0x073c
		"10100000",	-- 0x073d
		"11000110",	-- 0x073e
		"00001100",	-- 0x073f
		"10010010",	-- 0x0740
		"10100000",	-- 0x0741
		"00000000",	-- 0x0742
		"00000000",	-- 0x0743
		"00000000",	-- 0x0744
		"01010010",	-- 0x0745
		"01010011",	-- 0x0746
		"10011010",	-- 0x0747
		"00101100",	-- 0x0748
		"01110010",	-- 0x0749
		"10101101",	-- 0x074a
		"01110010",	-- 0x074b
		"00100011",	-- 0x074c
		"10000110",	-- 0x074d
		"00000001",	-- 0x074e
		"00000111",	-- 0x074f
		"10011010",	-- 0x0750
		"00000000",	-- 0x0751
		"10001011",	-- 0x0752
		"00000010",	-- 0x0753
		"11111111",	-- 0x0754
		"01110101",	-- 0x0755
		"01101011",	-- 0x0756
		"00110011",	-- 0x0757
		"00110000",	-- 0x0758
		"00000111",	-- 0x0759
		"00110011",	-- 0x075a
		"11110011",	-- 0x075b
		"00100111",	-- 0x075c
		"00000101",	-- 0x075d
		"11011011",	-- 0x075e
		"00101111",	-- 0x075f
		"11000011",	-- 0x0760
		"11001110",	-- 0x0761
		"11000111",	-- 0x0762
		"11001010",	-- 0x0763
		"11001010",	-- 0x0764
		"00010001",	-- 0x0765
		"10011010",	-- 0x0766
		"00101110",	-- 0x0767
		"11011010",	-- 0x0768
		"00100100",	-- 0x0769
		"11000010",	-- 0x076a
		"00111111",	-- 0x076b
		"11000110",	-- 0x076c
		"00011111",	-- 0x076d
		"10010010",	-- 0x076e
		"00100100",	-- 0x076f
		"11111010",	-- 0x0770
		"00000001",	-- 0x0771
		"11011101",	-- 0x0772
		"11000010",	-- 0x0773
		"11110100",	-- 0x0774
		"11000110",	-- 0x0775
		"01110100",	-- 0x0776
		"10110010",	-- 0x0777
		"00000001",	-- 0x0778
		"11011101",	-- 0x0779
		"10010010",	-- 0x077a
		"00010010",	-- 0x077b
		"11011010",	-- 0x077c
		"00000011",	-- 0x077d
		"11000010",	-- 0x077e
		"11111001",	-- 0x077f
		"11000110",	-- 0x0780
		"01111001",	-- 0x0781
		"10010010",	-- 0x0782
		"00000011",	-- 0x0783
		"00000111",	-- 0x0784
		"00110011",	-- 0x0785
		"11100011",	-- 0x0786
		"00010001",	-- 0x0787
		"00110011",	-- 0x0788
		"00011000",	-- 0x0789
		"00010000",	-- 0x078a
		"00110011",	-- 0x078b
		"11111100",	-- 0x078c
		"00010100",	-- 0x078d
		"00110011",	-- 0x078e
		"00110000",	-- 0x078f
		"00010011",	-- 0x0790
		"00110011",	-- 0x0791
		"00000000",	-- 0x0792
		"00011101",	-- 0x0793
		"10000110",	-- 0x0794
		"10000001",	-- 0x0795
		"11011110",	-- 0x0796
		"10011010",	-- 0x0797
		"00011000",	-- 0x0798
		"10000110",	-- 0x0799
		"10010010",	-- 0x079a
		"00000000",	-- 0x079b
		"10011010",	-- 0x079c
		"00011010",	-- 0x079d
		"00110101",	-- 0x079e
		"11110110",	-- 0x079f
		"00001100",	-- 0x07a0
		"00110111",	-- 0x07a1
		"00010000",	-- 0x07a2
		"00000110",	-- 0x07a3
		"00110111",	-- 0x07a4
		"00011001",	-- 0x07a5
		"00000011",	-- 0x07a6
		"00110101",	-- 0x07a7
		"00111001",	-- 0x07a8
		"00000011",	-- 0x07a9
		"01110111",	-- 0x07aa
		"01001011",	-- 0x07ab
		"10001100",	-- 0x07ac
		"01110101",	-- 0x07ad
		"01001011",	-- 0x07ae
		"01110001",	-- 0x07af
		"10101010",	-- 0x07b0
		"01000110",	-- 0x07b1
		"00000110",	-- 0x07b2
		"01110010",	-- 0x07b3
		"10111111",	-- 0x07b4
		"01110101",	-- 0x07b5
		"01000110",	-- 0x07b6
		"01110101",	-- 0x07b7
		"11010100",	-- 0x07b8
		"00110101",	-- 0x07b9
		"10101101",	-- 0x07ba
		"00000011",	-- 0x07bb
		"00110111",	-- 0x07bc
		"10101001",	-- 0x07bd
		"00000100",	-- 0x07be
		"01110101",	-- 0x07bf
		"10101101",	-- 0x07c0
		"01110010",	-- 0x07c1
		"10111110",	-- 0x07c2
		"00110111",	-- 0x07c3
		"00011001",	-- 0x07c4
		"00000010",	-- 0x07c5
		"01110010",	-- 0x07c6
		"11000000",	-- 0x07c7
		"00110101",	-- 0x07c8
		"10101010",	-- 0x07c9
		"00000011",	-- 0x07ca
		"00000011",	-- 0x07cb
		"11001000",	-- 0x07cc
		"01110011",	-- 0x07cd
		"01110001",	-- 0x07ce
		"11101010",	-- 0x07cf
		"01000111",	-- 0x07d0
		"00101101",	-- 0x07d1
		"01111001",	-- 0x07d2
		"01011010",	-- 0x07d3
		"10011100",	-- 0x07d4
		"01000110",	-- 0x07d5
		"00101000",	-- 0x07d6
		"10001111",	-- 0x07d7
		"00000011",	-- 0x07d8
		"00000000",	-- 0x07d9
		"10001101",	-- 0x07da
		"00000011",	-- 0x07db
		"00000100",	-- 0x07dc
		"01000100",	-- 0x07dd
		"00000111",	-- 0x07de
		"00011011",	-- 0x07df
		"00001000",	-- 0x07e0
		"01010110",	-- 0x07e1
		"01000111",	-- 0x07e2
		"11110110",	-- 0x07e3
		"01000000",	-- 0x07e4
		"00011001",	-- 0x07e5
		"10001111",	-- 0x07e6
		"00000000",	-- 0x07e7
		"10000000",	-- 0x07e8
		"10001101",	-- 0x07e9
		"00000000",	-- 0x07ea
		"10011110",	-- 0x07eb
		"01000100",	-- 0x07ec
		"00000111",	-- 0x07ed
		"00011011",	-- 0x07ee
		"00001000",	-- 0x07ef
		"01010110",	-- 0x07f0
		"01000111",	-- 0x07f1
		"11110110",	-- 0x07f2
		"01000000",	-- 0x07f3
		"00001010",	-- 0x07f4
		"11111011",	-- 0x07f5
		"00000011",	-- 0x07f6
		"00000000",	-- 0x07f7
		"10001111",	-- 0x07f8
		"11000011",	-- 0x07f9
		"11010011",	-- 0x07fa
		"00100001",	-- 0x07fb
		"10000100",	-- 0x07fc
		"01000100",	-- 0x07fd
		"00000010",	-- 0x07fe
		"01100001",	-- 0x07ff
		"00000111",	-- 0x0800
		"00110111",	-- 0x0801
		"10101010",	-- 0x0802
		"00000010",	-- 0x0803
		"01110111",	-- 0x0804
		"00010010",	-- 0x0805
		"01000000",	-- 0x0806
		"01101011",	-- 0x0807
		"01110010",	-- 0x0808
		"10011100",	-- 0x0809
		"10000110",	-- 0x080a
		"00000000",	-- 0x080b
		"11111111",	-- 0x080c
		"10001111",	-- 0x080d
		"00000000",	-- 0x080e
		"10000000",	-- 0x080f
		"10001010",	-- 0x0810
		"10001010",	-- 0x0811
		"10001010",	-- 0x0812
		"01110010",	-- 0x0813
		"01001011",	-- 0x0814
		"01110010",	-- 0x0815
		"01001100",	-- 0x0816
		"11011010",	-- 0x0817
		"10100000",	-- 0x0818
		"11000010",	-- 0x0819
		"00001100",	-- 0x081a
		"10010010",	-- 0x081b
		"10100000",	-- 0x081c
		"01110101",	-- 0x081d
		"10011101",	-- 0x081e
		"01110101",	-- 0x081f
		"01111000",	-- 0x0820
		"01110101",	-- 0x0821
		"00111101",	-- 0x0822
		"01110101",	-- 0x0823
		"10011000",	-- 0x0824
		"01110101",	-- 0x0825
		"10111000",	-- 0x0826
		"10000110",	-- 0x0827
		"10000000",	-- 0x0828
		"01111111",	-- 0x0829
		"10001111",	-- 0x082a
		"00000000",	-- 0x082b
		"10000110",	-- 0x082c
		"10001010",	-- 0x082d
		"10001101",	-- 0x082e
		"00000000",	-- 0x082f
		"10010100",	-- 0x0830
		"01000011",	-- 0x0831
		"11111010",	-- 0x0832
		"10000110",	-- 0x0833
		"00000000",	-- 0x0834
		"11111111",	-- 0x0835
		"10011010",	-- 0x0836
		"10010110",	-- 0x0837
		"10000110",	-- 0x0838
		"01100001",	-- 0x0839
		"10011110",	-- 0x083a
		"00110101",	-- 0x083b
		"00010000",	-- 0x083c
		"00000011",	-- 0x083d
		"10000110",	-- 0x083e
		"01010000",	-- 0x083f
		"10101111",	-- 0x0840
		"10011010",	-- 0x0841
		"10011000",	-- 0x0842
		"10000110",	-- 0x0843
		"01100110",	-- 0x0844
		"10011001",	-- 0x0845
		"10011010",	-- 0x0846
		"10011010",	-- 0x0847
		"10110010",	-- 0x0848
		"00000001",	-- 0x0849
		"10001110",	-- 0x084a
		"11011010",	-- 0x084b
		"10011110",	-- 0x084c
		"11000110",	-- 0x084d
		"00000001",	-- 0x084e
		"10010010",	-- 0x084f
		"10011110",	-- 0x0850
		"01010010",	-- 0x0851
		"10010010",	-- 0x0852
		"10011111",	-- 0x0853
		"10000110",	-- 0x0854
		"10101110",	-- 0x0855
		"01010001",	-- 0x0856
		"10111010",	-- 0x0857
		"00000011",	-- 0x0858
		"00000000",	-- 0x0859
		"10000110",	-- 0x085a
		"10101110",	-- 0x085b
		"01010001",	-- 0x085c
		"10111010",	-- 0x085d
		"00000011",	-- 0x085e
		"00000010",	-- 0x085f
		"00000101",	-- 0x0860
		"10000110",	-- 0x0861
		"10011010",	-- 0x0862
		"10011010",	-- 0x0863
		"10111010",	-- 0x0864
		"00000011",	-- 0x0865
		"00000100",	-- 0x0866
		"10110010",	-- 0x0867
		"00000011",	-- 0x0868
		"00000110",	-- 0x0869
		"00000111",	-- 0x086a
		"10000110",	-- 0x086b
		"01011010",	-- 0x086c
		"10100101",	-- 0x086d
		"10011010",	-- 0x086e
		"10011100",	-- 0x086f
		"01110101",	-- 0x0870
		"00010010",	-- 0x0871
		"01100011",	-- 0x0872
		"11111010",	-- 0x0873
		"00000001",	-- 0x0874
		"11011100",	-- 0x0875
		"01110001",	-- 0x0876
		"00010001",	-- 0x0877
		"01000110",	-- 0x0878
		"00000100",	-- 0x0879
		"11000110",	-- 0x087a
		"00000001",	-- 0x087b
		"01000000",	-- 0x087c
		"00000010",	-- 0x087d
		"11000010",	-- 0x087e
		"11111110",	-- 0x087f
		"10110010",	-- 0x0880
		"00000001",	-- 0x0881
		"11011100",	-- 0x0882
		"00000101",	-- 0x0883
		"01111001",	-- 0x0884
		"00111101",	-- 0x0885
		"11000111",	-- 0x0886
		"01000101",	-- 0x0887
		"00101011",	-- 0x0888
		"01010010",	-- 0x0889
		"01010011",	-- 0x088a
		"10011010",	-- 0x088b
		"01110100",	-- 0x088c
		"10011010",	-- 0x088d
		"11111000",	-- 0x088e
		"10111010",	-- 0x088f
		"00000001",	-- 0x0890
		"10100101",	-- 0x0891
		"00000001",	-- 0x0892
		"11110000",	-- 0x0893
		"00100000",	-- 0x0894
		"01110101",	-- 0x0895
		"00000110",	-- 0x0896
		"10000110",	-- 0x0897
		"00000000",	-- 0x0898
		"00000010",	-- 0x0899
		"10010111",	-- 0x089a
		"00000100",	-- 0x089b
		"10011010",	-- 0x089c
		"00001000",	-- 0x089d
		"01110101",	-- 0x089e
		"10000110",	-- 0x089f
		"01110101",	-- 0x08a0
		"10100110",	-- 0x08a1
		"01110101",	-- 0x08a2
		"11000110",	-- 0x08a3
		"01110101",	-- 0x08a4
		"11100110",	-- 0x08a5
		"01110010",	-- 0x08a6
		"00100001",	-- 0x08a7
		"01110101",	-- 0x08a8
		"10010011",	-- 0x08a9
		"01110101",	-- 0x08aa
		"10110100",	-- 0x08ab
		"00000111",	-- 0x08ac
		"01010010",	-- 0x08ad
		"01010011",	-- 0x08ae
		"10110010",	-- 0x08af
		"00000001",	-- 0x08b0
		"01101000",	-- 0x08b1
		"01000000",	-- 0x08b2
		"00000011",	-- 0x08b3
		"00000111",	-- 0x08b4
		"01100001",	-- 0x08b5
		"00001001",	-- 0x08b6
		"10011010",	-- 0x08b7
		"01011001",	-- 0x08b8
		"00000001",	-- 0x08b9
		"11000100",	-- 0x08ba
		"11011010",	-- 0x08bb
		"10010011",	-- 0x08bc
		"01011011",	-- 0x08bd
		"01000000",	-- 0x08be
		"00101110",	-- 0x08bf
		"10010110",	-- 0x08c0
		"11110110",	-- 0x08c1
		"11001100",	-- 0x08c2
		"00000011",	-- 0x08c3
		"01000100",	-- 0x08c4
		"00000011",	-- 0x08c5
		"10000110",	-- 0x08c6
		"00000011",	-- 0x08c7
		"00000000",	-- 0x08c8
		"10001110",	-- 0x08c9
		"11000100",	-- 0x08ca
		"11001010",	-- 0x08cb
		"01011000",	-- 0x08cc
		"01001011",	-- 0x08cd
		"00001101",	-- 0x08ce
		"00011100",	-- 0x08cf
		"00000110",	-- 0x08d0
		"01000000",	-- 0x08d1
		"11111001",	-- 0x08d2
		"10100100",	-- 0x08d3
		"10000100",	-- 0x08d4
		"01101010",	-- 0x08d5
		"01010101",	-- 0x08d6
		"01000011",	-- 0x08d7
		"00110100",	-- 0x08d8
		"00100111",	-- 0x08d9
		"00011100",	-- 0x08da
		"00010010",	-- 0x08db
		"00000001",	-- 0x08dc
		"11000100",	-- 0x08dd
		"11001100",	-- 0x08de
		"10001111",	-- 0x08df
		"11001000",	-- 0x08e0
		"11001001",	-- 0x08e1
		"01101110",	-- 0x08e2
		"00000001",	-- 0x08e3
		"11000100",	-- 0x08e4
		"01011001",	-- 0x08e5
		"00000100",	-- 0x08e6
		"11000000",	-- 0x08e7
		"01000000",	-- 0x08e8
		"01111110",	-- 0x08e9
		"00100001",	-- 0x08ea
		"00000000",	-- 0x08eb
		"00000110",	-- 0x08ec
		"01100011",	-- 0x08ed
		"11111010",	-- 0x08ee
		"00000001",	-- 0x08ef
		"11011100",	-- 0x08f0
		"11001110",	-- 0x08f1
		"00000001",	-- 0x08f2
		"01000110",	-- 0x08f3
		"00000010",	-- 0x08f4
		"01000000",	-- 0x08f5
		"00100001",	-- 0x08f6
		"10010110",	-- 0x08f7
		"01011001",	-- 0x08f8
		"10011110",	-- 0x08f9
		"01100000",	-- 0x08fa
		"01001010",	-- 0x08fb
		"00011001",	-- 0x08fc
		"11001100",	-- 0x08fd
		"00001001",	-- 0x08fe
		"01000101",	-- 0x08ff
		"00010101",	-- 0x0900
		"11001100",	-- 0x0901
		"00011001",	-- 0x0902
		"01000100",	-- 0x0903
		"00010001",	-- 0x0904
		"10011000",	-- 0x0905
		"01110100",	-- 0x0906
		"01000111",	-- 0x0907
		"00001111",	-- 0x0908
		"00010100",	-- 0x0909
		"00010101",	-- 0x090a
		"00000001",	-- 0x090b
		"11000100",	-- 0x090c
		"11010001",	-- 0x090d
		"10001001",	-- 0x090e
		"00000000",	-- 0x090f
		"00000000",	-- 0x0910
		"01000110",	-- 0x0911
		"00000001",	-- 0x0912
		"01010111",	-- 0x0913
		"10010111",	-- 0x0914
		"01110100",	-- 0x0915
		"10011010",	-- 0x0916
		"01110100",	-- 0x0917
		"01000000",	-- 0x0918
		"00100011",	-- 0x0919
		"01110101",	-- 0x091a
		"00011000",	-- 0x091b
		"10010110",	-- 0x091c
		"11111000",	-- 0x091d
		"10011000",	-- 0x091e
		"01011001",	-- 0x091f
		"01000100",	-- 0x0920
		"00000110",	-- 0x0921
		"01110111",	-- 0x0922
		"00011000",	-- 0x0923
		"01010100",	-- 0x0924
		"01010101",	-- 0x0925
		"10000100",	-- 0x0926
		"00000000",	-- 0x0927
		"00000001",	-- 0x0928
		"11000100",	-- 0x0929
		"11011101",	-- 0x092a
		"00010001",	-- 0x092b
		"00110111",	-- 0x092c
		"00011000",	-- 0x092d
		"00000001",	-- 0x092e
		"01010101",	-- 0x092f
		"11000001",	-- 0x0930
		"10000000",	-- 0x0931
		"10010011",	-- 0x0932
		"01011100",	-- 0x0933
		"10010110",	-- 0x0934
		"01011001",	-- 0x0935
		"10010111",	-- 0x0936
		"11111000",	-- 0x0937
		"00010100",	-- 0x0938
		"00010101",	-- 0x0939
		"10011010",	-- 0x093a
		"11111000",	-- 0x093b
		"01100011",	-- 0x093c
		"11011010",	-- 0x093d
		"01011011",	-- 0x093e
		"11001100",	-- 0x093f
		"00001000",	-- 0x0940
		"01000100",	-- 0x0941
		"00000010",	-- 0x0942
		"01110111",	-- 0x0943
		"00010110",	-- 0x0944
		"11001100",	-- 0x0945
		"00010000",	-- 0x0946
		"01000101",	-- 0x0947
		"00000010",	-- 0x0948
		"01110101",	-- 0x0949
		"00010110",	-- 0x094a
		"11001100",	-- 0x094b
		"00001100",	-- 0x094c
		"01000100",	-- 0x094d
		"00000010",	-- 0x094e
		"01110111",	-- 0x094f
		"10110000",	-- 0x0950
		"11001100",	-- 0x0951
		"00010100",	-- 0x0952
		"01000101",	-- 0x0953
		"00000010",	-- 0x0954
		"01110101",	-- 0x0955
		"10110000",	-- 0x0956
		"00110111",	-- 0x0957
		"00010110",	-- 0x0958
		"00000010",	-- 0x0959
		"01110010",	-- 0x095a
		"11010001",	-- 0x095b
		"11001100",	-- 0x095c
		"00001000",	-- 0x095d
		"01000101",	-- 0x095e
		"00000111",	-- 0x095f
		"00110101",	-- 0x0960
		"10110100",	-- 0x0961
		"00001000",	-- 0x0962
		"11001100",	-- 0x0963
		"00010000",	-- 0x0964
		"01000100",	-- 0x0965
		"00000100",	-- 0x0966
		"01110010",	-- 0x0967
		"11010000",	-- 0x0968
		"01110010",	-- 0x0969
		"11101010",	-- 0x096a
		"00110111",	-- 0x096b
		"01010110",	-- 0x096c
		"00000011",	-- 0x096d
		"01110111",	-- 0x096e
		"00010100",	-- 0x096f
		"10001100",	-- 0x0970
		"01110101",	-- 0x0971
		"00010100",	-- 0x0972
		"00110111",	-- 0x0973
		"00111001",	-- 0x0974
		"00011010",	-- 0x0975
		"11001010",	-- 0x0976
		"00011000",	-- 0x0977
		"01111001",	-- 0x0978
		"10010010",	-- 0x0979
		"01010111",	-- 0x097a
		"01000101",	-- 0x097b
		"00001000",	-- 0x097c
		"11011011",	-- 0x097d
		"01011011",	-- 0x097e
		"10001111",	-- 0x097f
		"11000010",	-- 0x0980
		"01010011",	-- 0x0981
		"00000001",	-- 0x0982
		"11000100",	-- 0x0983
		"01000111",	-- 0x0984
		"11011100",	-- 0x0985
		"10110001",	-- 0x0986
		"01000010",	-- 0x0987
		"00001001",	-- 0x0988
		"01110111",	-- 0x0989
		"01010110",	-- 0x098a
		"00110011",	-- 0x098b
		"11111110",	-- 0x098c
		"10110001",	-- 0x098d
		"01000000",	-- 0x098e
		"00000100",	-- 0x098f
		"01110010",	-- 0x0990
		"10110001",	-- 0x0991
		"01110101",	-- 0x0992
		"01010110",	-- 0x0993
		"01000000",	-- 0x0994
		"01000100",	-- 0x0995
		"00110111",	-- 0x0996
		"00111001",	-- 0x0997
		"00100100",	-- 0x0998
		"00110101",	-- 0x0999
		"10010111",	-- 0x099a
		"00100011",	-- 0x099b
		"00110101",	-- 0x099c
		"11110000",	-- 0x099d
		"00011011",	-- 0x099e
		"10110110",	-- 0x099f
		"00000001",	-- 0x09a0
		"01010000",	-- 0x09a1
		"00000001",	-- 0x09a2
		"11000100",	-- 0x09a3
		"11011011",	-- 0x09a4
		"01011010",	-- 0x09a5
		"11111011",	-- 0x09a6
		"00000001",	-- 0x09a7
		"00000001",	-- 0x09a8
		"00001001",	-- 0x09a9
		"01000011",	-- 0x09aa
		"00000010",	-- 0x09ab
		"01010111",	-- 0x09ac
		"01010000",	-- 0x09ad
		"00010100",	-- 0x09ae
		"00011000",	-- 0x09af
		"00001000",	-- 0x09b0
		"11001100",	-- 0x09b1
		"00010000",	-- 0x09b2
		"01000011",	-- 0x09b3
		"00000010",	-- 0x09b4
		"11001010",	-- 0x09b5
		"00010000",	-- 0x09b6
		"10110010",	-- 0x09b7
		"00000001",	-- 0x09b8
		"00000001",	-- 0x09b9
		"01110111",	-- 0x09ba
		"10010111",	-- 0x09bb
		"10001100",	-- 0x09bc
		"01110101",	-- 0x09bd
		"10010111",	-- 0x09be
		"11111011",	-- 0x09bf
		"00000001",	-- 0x09c0
		"00000001",	-- 0x09c1
		"00010001",	-- 0x09c2
		"11001101",	-- 0x09c3
		"00000100",	-- 0x09c4
		"01000100",	-- 0x09c5
		"00000010",	-- 0x09c6
		"11001011",	-- 0x09c7
		"00000100",	-- 0x09c8
		"00010001",	-- 0x09c9
		"00010001",	-- 0x09ca
		"11111101",	-- 0x09cb
		"00000001",	-- 0x09cc
		"01010000",	-- 0x09cd
		"01000010",	-- 0x09ce
		"00000111",	-- 0x09cf
		"01110001",	-- 0x09d0
		"10010000",	-- 0x09d1
		"01000111",	-- 0x09d2
		"00000101",	-- 0x09d3
		"01110010",	-- 0x09d4
		"10110001",	-- 0x09d5
		"10001100",	-- 0x09d6
		"01110101",	-- 0x09d7
		"10010000",	-- 0x09d8
		"01100011",	-- 0x09d9
		"00110101",	-- 0x09da
		"01011001",	-- 0x09db
		"00000010",	-- 0x09dc
		"01110010",	-- 0x09dd
		"10111000",	-- 0x09de
		"01111001",	-- 0x09df
		"00110001",	-- 0x09e0
		"10111000",	-- 0x09e1
		"01000101",	-- 0x09e2
		"00000011",	-- 0x09e3
		"01110111",	-- 0x09e4
		"11010101",	-- 0x09e5
		"10001100",	-- 0x09e6
		"01110101",	-- 0x09e7
		"11010101",	-- 0x09e8
		"00110101",	-- 0x09e9
		"11010101",	-- 0x09ea
		"00000010",	-- 0x09eb
		"01110010",	-- 0x09ec
		"10111001",	-- 0x09ed
		"11111010",	-- 0x09ee
		"00000001",	-- 0x09ef
		"11010111",	-- 0x09f0
		"10010010",	-- 0x09f1
		"01001110",	-- 0x09f2
		"00110101",	-- 0x09f3
		"01111001",	-- 0x09f4
		"00000100",	-- 0x09f5
		"01110010",	-- 0x09f6
		"10101111",	-- 0x09f7
		"01000000",	-- 0x09f8
		"00000101",	-- 0x09f9
		"01111001",	-- 0x09fa
		"01011100",	-- 0x09fb
		"11010000",	-- 0x09fc
		"01000100",	-- 0x09fd
		"00000101",	-- 0x09fe
		"00110111",	-- 0x09ff
		"11010110",	-- 0x0a00
		"00011001",	-- 0x0a01
		"01000000",	-- 0x0a02
		"00001101",	-- 0x0a03
		"00110101",	-- 0x0a04
		"11010110",	-- 0x0a05
		"00010010",	-- 0x0a06
		"01111001",	-- 0x0a07
		"00110001",	-- 0x0a08
		"10101111",	-- 0x0a09
		"01000101",	-- 0x0a0a
		"00001111",	-- 0x0a0b
		"01111001",	-- 0x0a0c
		"01011100",	-- 0x0a0d
		"11010000",	-- 0x0a0e
		"01000101",	-- 0x0a0f
		"00001010",	-- 0x0a10
		"01110001",	-- 0x0a11
		"11010110",	-- 0x0a12
		"01000111",	-- 0x0a13
		"00000010",	-- 0x0a14
		"01110101",	-- 0x0a15
		"11010110",	-- 0x0a16
		"01110111",	-- 0x0a17
		"11111110",	-- 0x0a18
		"01110010",	-- 0x0a19
		"10101111",	-- 0x0a1a
		"01110101",	-- 0x0a1b
		"11010000",	-- 0x0a1c
		"01110111",	-- 0x0a1d
		"11010010",	-- 0x0a1e
		"01110101",	-- 0x0a1f
		"00111110",	-- 0x0a20
		"11011010",	-- 0x0a21
		"01001110",	-- 0x0a22
		"10110010",	-- 0x0a23
		"00000001",	-- 0x0a24
		"11010111",	-- 0x0a25
		"00000001",	-- 0x0a26
		"11100100",	-- 0x0a27
		"01010100",	-- 0x0a28
		"00000001",	-- 0x0a29
		"11100101",	-- 0x0a2a
		"01010001",	-- 0x0a2b
		"00000001",	-- 0x0a2c
		"11111100",	-- 0x0a2d
		"00111000",	-- 0x0a2e
		"00000001",	-- 0x0a2f
		"11010010",	-- 0x0a30
		"11000101",	-- 0x0a31
		"11111010",	-- 0x0a32
		"00000001",	-- 0x0a33
		"11010101",	-- 0x0a34
		"10010010",	-- 0x0a35
		"01001110",	-- 0x0a36
		"00110111",	-- 0x0a37
		"00010011",	-- 0x0a38
		"00000011",	-- 0x0a39
		"01110111",	-- 0x0a3a
		"01110100",	-- 0x0a3b
		"10001100",	-- 0x0a3c
		"01110101",	-- 0x0a3d
		"01110100",	-- 0x0a3e
		"01110101",	-- 0x0a3f
		"10111110",	-- 0x0a40
		"01110101",	-- 0x0a41
		"00011110",	-- 0x0a42
		"11001011",	-- 0x0a43
		"00001100",	-- 0x0a44
		"01111001",	-- 0x0a45
		"01011100",	-- 0x0a46
		"11010000",	-- 0x0a47
		"01000100",	-- 0x0a48
		"00010010",	-- 0x0a49
		"00110111",	-- 0x0a4a
		"01010110",	-- 0x0a4b
		"00010111",	-- 0x0a4c
		"01111001",	-- 0x0a4d
		"11100001",	-- 0x0a4e
		"01010111",	-- 0x0a4f
		"01000101",	-- 0x0a50
		"00010010",	-- 0x0a51
		"01111001",	-- 0x0a52
		"00000010",	-- 0x0a53
		"01011101",	-- 0x0a54
		"01000010",	-- 0x0a55
		"00001101",	-- 0x0a56
		"01010011",	-- 0x0a57
		"01110111",	-- 0x0a58
		"00011110",	-- 0x0a59
		"01000000",	-- 0x0a5a
		"00001000",	-- 0x0a5b
		"00110101",	-- 0x0a5c
		"00010011",	-- 0x0a5d
		"00000011",	-- 0x0a5e
		"00110101",	-- 0x0a5f
		"00010100",	-- 0x0a60
		"00000010",	-- 0x0a61
		"11001011",	-- 0x0a62
		"00001100",	-- 0x0a63
		"11111010",	-- 0x0a64
		"00000001",	-- 0x0a65
		"01001000",	-- 0x0a66
		"00110101",	-- 0x0a67
		"00011110",	-- 0x0a68
		"00001000",	-- 0x0a69
		"01111001",	-- 0x0a6a
		"00011001",	-- 0x0a6b
		"01011101",	-- 0x0a6c
		"01000100",	-- 0x0a6d
		"00001001",	-- 0x0a6e
		"00110101",	-- 0x0a6f
		"10011001",	-- 0x0a70
		"00000110",	-- 0x0a71
		"11001100",	-- 0x0a72
		"01000100",	-- 0x0a73
		"01000100",	-- 0x0a74
		"00000010",	-- 0x0a75
		"11001010",	-- 0x0a76
		"01000100",	-- 0x0a77
		"00110101",	-- 0x0a78
		"00010011",	-- 0x0a79
		"00101111",	-- 0x0a7a
		"00001000",	-- 0x0a7b
		"11001011",	-- 0x0a7c
		"01000100",	-- 0x0a7d
		"00110101",	-- 0x0a7e
		"00011110",	-- 0x0a7f
		"00010010",	-- 0x0a80
		"11001011",	-- 0x0a81
		"01010000",	-- 0x0a82
		"01111001",	-- 0x0a83
		"00010001",	-- 0x0a84
		"01011101",	-- 0x0a85
		"01000101",	-- 0x0a86
		"00001011",	-- 0x0a87
		"01111001",	-- 0x0a88
		"00011110",	-- 0x0a89
		"01011101",	-- 0x0a8a
		"01000100",	-- 0x0a8b
		"00001010",	-- 0x0a8c
		"00110101",	-- 0x0a8d
		"11010110",	-- 0x0a8e
		"00000011",	-- 0x0a8f
		"00110101",	-- 0x0a90
		"10011001",	-- 0x0a91
		"00000100",	-- 0x0a92
		"00001011",	-- 0x0a93
		"01000100",	-- 0x0a94
		"00000001",	-- 0x0a95
		"01011010",	-- 0x0a96
		"00110111",	-- 0x0a97
		"01010110",	-- 0x0a98
		"00111010",	-- 0x0a99
		"11011100",	-- 0x0a9a
		"01011011",	-- 0x0a9b
		"01000010",	-- 0x0a9c
		"00110110",	-- 0x0a9d
		"01111001",	-- 0x0a9e
		"00011000",	-- 0x0a9f
		"10110110",	-- 0x0aa0
		"01000101",	-- 0x0aa1
		"00110001",	-- 0x0aa2
		"01111001",	-- 0x0aa3
		"00011000",	-- 0x0aa4
		"10110111",	-- 0x0aa5
		"01000101",	-- 0x0aa6
		"00101100",	-- 0x0aa7
		"01000000",	-- 0x0aa8
		"00110011",	-- 0x0aa9
		"00110111",	-- 0x0aaa
		"01010110",	-- 0x0aab
		"00100111",	-- 0x0aac
		"01111001",	-- 0x0aad
		"00011000",	-- 0x0aae
		"10110110",	-- 0x0aaf
		"01000101",	-- 0x0ab0
		"00100010",	-- 0x0ab1
		"01111001",	-- 0x0ab2
		"00011000",	-- 0x0ab3
		"10110111",	-- 0x0ab4
		"01000101",	-- 0x0ab5
		"00011101",	-- 0x0ab6
		"11011100",	-- 0x0ab7
		"01011011",	-- 0x0ab8
		"01000011",	-- 0x0ab9
		"00000111",	-- 0x0aba
		"01110111",	-- 0x0abb
		"10111110",	-- 0x0abc
		"00110011",	-- 0x0abd
		"01100110",	-- 0x0abe
		"01100000",	-- 0x0abf
		"01000000",	-- 0x0ac0
		"00010010",	-- 0x0ac1
		"01111001",	-- 0x0ac2
		"00101100",	-- 0x0ac3
		"01011011",	-- 0x0ac4
		"01000100",	-- 0x0ac5
		"00010110",	-- 0x0ac6
		"01111001",	-- 0x0ac7
		"00100011",	-- 0x0ac8
		"01011101",	-- 0x0ac9
		"01000100",	-- 0x0aca
		"00010001",	-- 0x0acb
		"01111001",	-- 0x0acc
		"10001011",	-- 0x0acd
		"01011100",	-- 0x0ace
		"01000101",	-- 0x0acf
		"00001100",	-- 0x0ad0
		"00000001",	-- 0x0ad1
		"11001101",	-- 0x0ad2
		"10111001",	-- 0x0ad3
		"00000001",	-- 0x0ad4
		"11001101",	-- 0x0ad5
		"01101000",	-- 0x0ad6
		"01110010",	-- 0x0ad7
		"11001110",	-- 0x0ad8
		"01110101",	-- 0x0ad9
		"00010011",	-- 0x0ada
		"01000000",	-- 0x0adb
		"00000101",	-- 0x0adc
		"01110111",	-- 0x0add
		"00010011",	-- 0x0ade
		"00110011",	-- 0x0adf
		"10000000",	-- 0x0ae0
		"01100000",	-- 0x0ae1
		"11011010",	-- 0x0ae2
		"01100000",	-- 0x0ae3
		"01001011",	-- 0x0ae4
		"00010101",	-- 0x0ae5
		"00110111",	-- 0x0ae6
		"01010110",	-- 0x0ae7
		"00010010",	-- 0x0ae8
		"01111001",	-- 0x0ae9
		"11011100",	-- 0x0aea
		"01010111",	-- 0x0aeb
		"01000101",	-- 0x0aec
		"00001101",	-- 0x0aed
		"01111001",	-- 0x0aee
		"00000101",	-- 0x0aef
		"01011101",	-- 0x0af0
		"01000101",	-- 0x0af1
		"00001000",	-- 0x0af2
		"01111001",	-- 0x0af3
		"10000111",	-- 0x0af4
		"01011100",	-- 0x0af5
		"01000011",	-- 0x0af6
		"00000110",	-- 0x0af7
		"00000001",	-- 0x0af8
		"11001101",	-- 0x0af9
		"10111110",	-- 0x0afa
		"00110011",	-- 0x0afb
		"10000000",	-- 0x0afc
		"01100000",	-- 0x0afd
		"01000000",	-- 0x0afe
		"00011110",	-- 0x0aff
		"11011010",	-- 0x0b00
		"01100000",	-- 0x0b01
		"11000000",	-- 0x0b02
		"00000010",	-- 0x0b03
		"01001010",	-- 0x0b04
		"00000010",	-- 0x0b05
		"11001010",	-- 0x0b06
		"10000000",	-- 0x0b07
		"10010010",	-- 0x0b08
		"01100000",	-- 0x0b09
		"01100011",	-- 0x0b0a
		"10001111",	-- 0x0b0b
		"11000001",	-- 0x0b0c
		"01000111",	-- 0x0b0d
		"00000001",	-- 0x0b0e
		"11000100",	-- 0x0b0f
		"00111100",	-- 0x0b10
		"00110111",	-- 0x0b11
		"11010110",	-- 0x0b12
		"00000110",	-- 0x0b13
		"11001100",	-- 0x0b14
		"00111100",	-- 0x0b15
		"01000100",	-- 0x0b16
		"00000010",	-- 0x0b17
		"11001010",	-- 0x0b18
		"00111100",	-- 0x0b19
		"10110010",	-- 0x0b1a
		"00000001",	-- 0x0b1b
		"01001000",	-- 0x0b1c
		"01100011",	-- 0x0b1d
		"00000001",	-- 0x0b1e
		"11101111",	-- 0x0b1f
		"00101100",	-- 0x0b20
		"10110110",	-- 0x0b21
		"00000001",	-- 0x0b22
		"00001010",	-- 0x0b23
		"10001001",	-- 0x0b24
		"00000000",	-- 0x0b25
		"10101111",	-- 0x0b26
		"01000011",	-- 0x0b27
		"00000010",	-- 0x0b28
		"01110010",	-- 0x0b29
		"11010110",	-- 0x0b2a
		"11001010",	-- 0x0b2b
		"01100000",	-- 0x0b2c
		"00110111",	-- 0x0b2d
		"00110011",	-- 0x0b2e
		"00000010",	-- 0x0b2f
		"11001010",	-- 0x0b30
		"01011100",	-- 0x0b31
		"11011100",	-- 0x0b32
		"01011011",	-- 0x0b33
		"01000010",	-- 0x0b34
		"00001111",	-- 0x0b35
		"11011010",	-- 0x0b36
		"01100000",	-- 0x0b37
		"01001010",	-- 0x0b38
		"00001011",	-- 0x0b39
		"00110101",	-- 0x0b3a
		"00010011",	-- 0x0b3b
		"00001000",	-- 0x0b3c
		"10111110",	-- 0x0b3d
		"00000001",	-- 0x0b3e
		"00001010",	-- 0x0b3f
		"10001100",	-- 0x0b40
		"00000001",	-- 0x0b41
		"00100000",	-- 0x0b42
		"01000101",	-- 0x0b43
		"00001000",	-- 0x0b44
		"01110010",	-- 0x0b45
		"11101011",	-- 0x0b46
		"01110101",	-- 0x0b47
		"00111110",	-- 0x0b48
		"01110101",	-- 0x0b49
		"00110011",	-- 0x0b4a
		"01000000",	-- 0x0b4b
		"00111101",	-- 0x0b4c
		"10001100",	-- 0x0b4d
		"00000000",	-- 0x0b4e
		"11100001",	-- 0x0b4f
		"01000100",	-- 0x0b50
		"00000010",	-- 0x0b51
		"01110111",	-- 0x0b52
		"00111110",	-- 0x0b53
		"10001100",	-- 0x0b54
		"00000001",	-- 0x0b55
		"00100000",	-- 0x0b56
		"01000101",	-- 0x0b57
		"00000010",	-- 0x0b58
		"01110101",	-- 0x0b59
		"00111110",	-- 0x0b5a
		"01111001",	-- 0x0b5b
		"00001010",	-- 0x0b5c
		"01011101",	-- 0x0b5d
		"01000101",	-- 0x0b5e
		"00000011",	-- 0x0b5f
		"00110101",	-- 0x0b60
		"00111110",	-- 0x0b61
		"00000010",	-- 0x0b62
		"01110010",	-- 0x0b63
		"11101011",	-- 0x0b64
		"01111001",	-- 0x0b65
		"00011000",	-- 0x0b66
		"10110110",	-- 0x0b67
		"01000101",	-- 0x0b68
		"11011111",	-- 0x0b69
		"01111001",	-- 0x0b6a
		"00011000",	-- 0x0b6b
		"10110111",	-- 0x0b6c
		"01000101",	-- 0x0b6d
		"11011010",	-- 0x0b6e
		"11011011",	-- 0x0b6f
		"01011011",	-- 0x0b70
		"10001111",	-- 0x0b71
		"11000001",	-- 0x0b72
		"01001101",	-- 0x0b73
		"00000001",	-- 0x0b74
		"11000100",	-- 0x0b75
		"01000100",	-- 0x0b76
		"11011100",	-- 0x0b77
		"11010110",	-- 0x0b78
		"01000011",	-- 0x0b79
		"00001101",	-- 0x0b7a
		"11001010",	-- 0x0b7b
		"00000101",	-- 0x0b7c
		"01111001",	-- 0x0b7d
		"01111000",	-- 0x0b7e
		"01011011",	-- 0x0b7f
		"01000100",	-- 0x0b80
		"00000010",	-- 0x0b81
		"11001010",	-- 0x0b82
		"00010100",	-- 0x0b83
		"11011100",	-- 0x0b84
		"11101011",	-- 0x0b85
		"01000010",	-- 0x0b86
		"00000010",	-- 0x0b87
		"01110111",	-- 0x0b88
		"00110011",	-- 0x0b89
		"01111001",	-- 0x0b8a
		"00001010",	-- 0x0b8b
		"01011101",	-- 0x0b8c
		"01000100",	-- 0x0b8d
		"00000110",	-- 0x0b8e
		"01111001",	-- 0x0b8f
		"00111100",	-- 0x0b90
		"01011011",	-- 0x0b91
		"01000100",	-- 0x0b92
		"00000101",	-- 0x0b93
		"10001100",	-- 0x0b94
		"01110101",	-- 0x0b95
		"01111110",	-- 0x0b96
		"01110101",	-- 0x0b97
		"10011110",	-- 0x0b98
		"00110101",	-- 0x0b99
		"11010011",	-- 0x0b9a
		"00100001",	-- 0x0b9b
		"01111001",	-- 0x0b9c
		"11011100",	-- 0x0b9d
		"01010111",	-- 0x0b9e
		"01000101",	-- 0x0b9f
		"00011100",	-- 0x0ba0
		"01111001",	-- 0x0ba1
		"00000000",	-- 0x0ba2
		"01011101",	-- 0x0ba3
		"01000110",	-- 0x0ba4
		"00010111",	-- 0x0ba5
		"00110101",	-- 0x0ba6
		"01111011",	-- 0x0ba7
		"00010100",	-- 0x0ba8
		"11011011",	-- 0x0ba9
		"01011001",	-- 0x0baa
		"11001101",	-- 0x0bab
		"00011000",	-- 0x0bac
		"01000101",	-- 0x0bad
		"00001110",	-- 0x0bae
		"11001101",	-- 0x0baf
		"01100100",	-- 0x0bb0
		"01000100",	-- 0x0bb1
		"00001010",	-- 0x0bb2
		"10001111",	-- 0x0bb3
		"11000001",	-- 0x0bb4
		"11100001",	-- 0x0bb5
		"00000001",	-- 0x0bb6
		"11000100",	-- 0x0bb7
		"01000100",	-- 0x0bb8
		"11011100",	-- 0x0bb9
		"01010000",	-- 0x0bba
		"01000011",	-- 0x0bbb
		"00000100",	-- 0x0bbc
		"01110010",	-- 0x0bbd
		"11001111",	-- 0x0bbe
		"01000000",	-- 0x0bbf
		"00001001",	-- 0x0bc0
		"01111001",	-- 0x0bc1
		"11110100",	-- 0x0bc2
		"11001111",	-- 0x0bc3
		"01000101",	-- 0x0bc4
		"00000100",	-- 0x0bc5
		"01110111",	-- 0x0bc6
		"10011110",	-- 0x0bc7
		"01110111",	-- 0x0bc8
		"01111110",	-- 0x0bc9
		"00110101",	-- 0x0bca
		"00010000",	-- 0x0bcb
		"00100010",	-- 0x0bcc
		"10000110",	-- 0x0bcd
		"00111100",	-- 0x0bce
		"01000110",	-- 0x0bcf
		"10011110",	-- 0x0bd0
		"01010111",	-- 0x0bd1
		"10001100",	-- 0x0bd2
		"11110011",	-- 0x0bd3
		"00000000",	-- 0x0bd4
		"01000101",	-- 0x0bd5
		"00000011",	-- 0x0bd6
		"10000110",	-- 0x0bd7
		"00101000",	-- 0x0bd8
		"00110010",	-- 0x0bd9
		"10011010",	-- 0x0bda
		"01111000",	-- 0x0bdb
		"01111001",	-- 0x0bdc
		"11011100",	-- 0x0bdd
		"01010111",	-- 0x0bde
		"01000101",	-- 0x0bdf
		"00001110",	-- 0x0be0
		"00110101",	-- 0x0be1
		"01010110",	-- 0x0be2
		"00001011",	-- 0x0be3
		"01111001",	-- 0x0be4
		"00001010",	-- 0x0be5
		"01011101",	-- 0x0be6
		"01000100",	-- 0x0be7
		"00000110",	-- 0x0be8
		"00110101",	-- 0x0be9
		"10011110",	-- 0x0bea
		"00000011",	-- 0x0beb
		"00110101",	-- 0x0bec
		"11010010",	-- 0x0bed
		"00001000",	-- 0x0bee
		"01010010",	-- 0x0bef
		"10010010",	-- 0x0bf0
		"01101000",	-- 0x0bf1
		"00000001",	-- 0x0bf2
		"11001100",	-- 0x0bf3
		"10010011",	-- 0x0bf4
		"01000000",	-- 0x0bf5
		"00110110",	-- 0x0bf6
		"11011011",	-- 0x0bf7
		"01011001",	-- 0x0bf8
		"11011010",	-- 0x0bf9
		"01101000",	-- 0x0bfa
		"11001100",	-- 0x0bfb
		"11111111",	-- 0x0bfc
		"01000100",	-- 0x0bfd
		"00001010",	-- 0x0bfe
		"11001010",	-- 0x0bff
		"10010100",	-- 0x0c00
		"00001011",	-- 0x0c01
		"01000011",	-- 0x0c02
		"00001101",	-- 0x0c03
		"00110111",	-- 0x0c04
		"11010011",	-- 0x0c05
		"11101011",	-- 0x0c06
		"01000000",	-- 0x0c07
		"00010010",	-- 0x0c08
		"11011010",	-- 0x0c09
		"11111000",	-- 0x0c0a
		"11011101",	-- 0x0c0b
		"01111001",	-- 0x0c0c
		"01000101",	-- 0x0c0d
		"00000010",	-- 0x0c0e
		"01110111",	-- 0x0c0f
		"01011110",	-- 0x0c10
		"01110001",	-- 0x0c11
		"11010011",	-- 0x0c12
		"01000110",	-- 0x0c13
		"00000110",	-- 0x0c14
		"01110010",	-- 0x0c15
		"11001101",	-- 0x0c16
		"11001011",	-- 0x0c17
		"00000000",	-- 0x0c18
		"01000000",	-- 0x0c19
		"00000011",	-- 0x0c1a
		"10110110",	-- 0x0c1b
		"00000001",	-- 0x0c1c
		"01001001",	-- 0x0c1d
		"11011100",	-- 0x0c1e
		"01111000",	-- 0x0c1f
		"01000100",	-- 0x0c20
		"00000010",	-- 0x0c21
		"11011010",	-- 0x0c22
		"01111000",	-- 0x0c23
		"11001101",	-- 0x0c24
		"00011110",	-- 0x0c25
		"01000011",	-- 0x0c26
		"00000010",	-- 0x0c27
		"11001011",	-- 0x0c28
		"00011110",	-- 0x0c29
		"10111010",	-- 0x0c2a
		"00000001",	-- 0x0c2b
		"01001001",	-- 0x0c2c
		"00110111",	-- 0x0c2d
		"01010011",	-- 0x0c2e
		"00001001",	-- 0x0c2f
		"11110100",	-- 0x0c30
		"00000001",	-- 0x0c31
		"01001010",	-- 0x0c32
		"11001100",	-- 0x0c33
		"00011110",	-- 0x0c34
		"01000100",	-- 0x0c35
		"00000010",	-- 0x0c36
		"11001010",	-- 0x0c37
		"00011110",	-- 0x0c38
		"11011100",	-- 0x0c39
		"01011001",	-- 0x0c3a
		"01000010",	-- 0x0c3b
		"00000101",	-- 0x0c3c
		"01110111",	-- 0x0c3d
		"01010011",	-- 0x0c3e
		"01110111",	-- 0x0c3f
		"01011110",	-- 0x0c40
		"10001100",	-- 0x0c41
		"01110101",	-- 0x0c42
		"01010011",	-- 0x0c43
		"01111001",	-- 0x0c44
		"00111101",	-- 0x0c45
		"11001101",	-- 0x0c46
		"01000101",	-- 0x0c47
		"01001000",	-- 0x0c48
		"01110010",	-- 0x0c49
		"11001101",	-- 0x0c4a
		"00110111",	-- 0x0c4b
		"01011110",	-- 0x0c4c
		"00010111",	-- 0x0c4d
		"00110111",	-- 0x0c4e
		"11010011",	-- 0x0c4f
		"00010111",	-- 0x0c50
		"10110110",	-- 0x0c51
		"00000001",	-- 0x0c52
		"01001001",	-- 0x0c53
		"11000100",	-- 0x0c54
		"00000001",	-- 0x0c55
		"01000100",	-- 0x0c56
		"00000010",	-- 0x0c57
		"11011010",	-- 0x0c58
		"01111000",	-- 0x0c59
		"11000001",	-- 0x0c5a
		"00000001",	-- 0x0c5b
		"01000100",	-- 0x0c5c
		"00000010",	-- 0x0c5d
		"11001011",	-- 0x0c5e
		"00011110",	-- 0x0c5f
		"10111010",	-- 0x0c60
		"00000001",	-- 0x0c61
		"01001001",	-- 0x0c62
		"01000000",	-- 0x0c63
		"00101010",	-- 0x0c64
		"00000001",	-- 0x0c65
		"11001100",	-- 0x0c66
		"10010011",	-- 0x0c67
		"11011010",	-- 0x0c68
		"01111001",	-- 0x0c69
		"11011100",	-- 0x0c6a
		"01011001",	-- 0x0c6b
		"01000011",	-- 0x0c6c
		"00000111",	-- 0x0c6d
		"11011010",	-- 0x0c6e
		"01101000",	-- 0x0c6f
		"01000111",	-- 0x0c70
		"00000001",	-- 0x0c71
		"01010000",	-- 0x0c72
		"01000000",	-- 0x0c73
		"00011000",	-- 0x0c74
		"10001111",	-- 0x0c75
		"11000001",	-- 0x0c76
		"11100111",	-- 0x0c77
		"11011011",	-- 0x0c78
		"01011001",	-- 0x0c79
		"00000001",	-- 0x0c7a
		"11000100",	-- 0x0c7b
		"01000111",	-- 0x0c7c
		"10011110",	-- 0x0c7d
		"01010111",	-- 0x0c7e
		"10001100",	-- 0x0c7f
		"11110101",	-- 0x0c80
		"11000000",	-- 0x0c81
		"01000101",	-- 0x0c82
		"00000011",	-- 0x0c83
		"00010010",	-- 0x0c84
		"01000101",	-- 0x0c85
		"00000100",	-- 0x0c86
		"11010000",	-- 0x0c87
		"01101000",	-- 0x0c88
		"01000100",	-- 0x0c89
		"00000010",	-- 0x0c8a
		"11001010",	-- 0x0c8b
		"11111111",	-- 0x0c8c
		"10010010",	-- 0x0c8d
		"01101000",	-- 0x0c8e
		"01110101",	-- 0x0c8f
		"01011110",	-- 0x0c90
		"01000000",	-- 0x0c91
		"00001001",	-- 0x0c92
		"01110101",	-- 0x0c93
		"11010011",	-- 0x0c94
		"10000110",	-- 0x0c95
		"10010100",	-- 0x0c96
		"00000000",	-- 0x0c97
		"10111010",	-- 0x0c98
		"00000001",	-- 0x0c99
		"01001001",	-- 0x0c9a
		"01100011",	-- 0x0c9b
		"00000001",	-- 0x0c9c
		"11101110",	-- 0x0c9d
		"10101000",	-- 0x0c9e
		"00110111",	-- 0x0c9f
		"01110011",	-- 0x0ca0
		"00010001",	-- 0x0ca1
		"01111001",	-- 0x0ca2
		"10110100",	-- 0x0ca3
		"01011101",	-- 0x0ca4
		"01000100",	-- 0x0ca5
		"00000101",	-- 0x0ca6
		"01111001",	-- 0x0ca7
		"00001000",	-- 0x0ca8
		"11100001",	-- 0x0ca9
		"01000100",	-- 0x0caa
		"00000101",	-- 0x0cab
		"01111001",	-- 0x0cac
		"00101000",	-- 0x0cad
		"01011001",	-- 0x0cae
		"01000100",	-- 0x0caf
		"00000100",	-- 0x0cb0
		"01110101",	-- 0x0cb1
		"01110011",	-- 0x0cb2
		"01110010",	-- 0x0cb3
		"11100001",	-- 0x0cb4
		"01000000",	-- 0x0cb5
		"00011010",	-- 0x0cb6
		"01010010",	-- 0x0cb7
		"01111001",	-- 0x0cb8
		"10110100",	-- 0x0cb9
		"01011101",	-- 0x0cba
		"01000101",	-- 0x0cbb
		"00000110",	-- 0x0cbc
		"11011010",	-- 0x0cbd
		"01101110",	-- 0x0cbe
		"01010110",	-- 0x0cbf
		"01000110",	-- 0x0cc0
		"00000001",	-- 0x0cc1
		"01010000",	-- 0x0cc2
		"10010010",	-- 0x0cc3
		"01101110",	-- 0x0cc4
		"11001100",	-- 0x0cc5
		"00000110",	-- 0x0cc6
		"01000101",	-- 0x0cc7
		"00000111",	-- 0x0cc8
		"01111001",	-- 0x0cc9
		"01010000",	-- 0x0cca
		"01011001",	-- 0x0ccb
		"01000101",	-- 0x0ccc
		"00000010",	-- 0x0ccd
		"01110111",	-- 0x0cce
		"01110011",	-- 0x0ccf
		"01100011",	-- 0x0cd0
		"00000001",	-- 0x0cd1
		"11101110",	-- 0x0cd2
		"10010011",	-- 0x0cd3
		"01000000",	-- 0x0cd4
		"00100101",	-- 0x0cd5
		"10001111",	-- 0x0cd6
		"11000001",	-- 0x0cd7
		"11101111",	-- 0x0cd8
		"10010110",	-- 0x0cd9
		"01011001",	-- 0x0cda
		"00000001",	-- 0x0cdb
		"11000100",	-- 0x0cdc
		"00101111",	-- 0x0cdd
		"00110111",	-- 0x0cde
		"11110011",	-- 0x0cdf
		"00000010",	-- 0x0ce0
		"11000100",	-- 0x0ce1
		"00001101",	-- 0x0ce2
		"11011100",	-- 0x0ce3
		"01010000",	-- 0x0ce4
		"01000011",	-- 0x0ce5
		"00000010",	-- 0x0ce6
		"01110010",	-- 0x0ce7
		"10111100",	-- 0x0ce8
		"10001111",	-- 0x0ce9
		"11000001",	-- 0x0cea
		"11110101",	-- 0x0ceb
		"10010110",	-- 0x0cec
		"01011001",	-- 0x0ced
		"00000001",	-- 0x0cee
		"11000100",	-- 0x0cef
		"00101111",	-- 0x0cf0
		"11011100",	-- 0x0cf1
		"10111100",	-- 0x0cf2
		"01000010",	-- 0x0cf3
		"00000011",	-- 0x0cf4
		"01110111",	-- 0x0cf5
		"11110011",	-- 0x0cf6
		"10001100",	-- 0x0cf7
		"01110101",	-- 0x0cf8
		"11110011",	-- 0x0cf9
		"01100011",	-- 0x0cfa
		"00110111",	-- 0x0cfb
		"11110011",	-- 0x0cfc
		"00001001",	-- 0x0cfd
		"01111001",	-- 0x0cfe
		"00011000",	-- 0x0cff
		"11000011",	-- 0x0d00
		"01000101",	-- 0x0d01
		"00000110",	-- 0x0d02
		"01110111",	-- 0x0d03
		"11111110",	-- 0x0d04
		"01000000",	-- 0x0d05
		"00000100",	-- 0x0d06
		"01110010",	-- 0x0d07
		"11000011",	-- 0x0d08
		"01110101",	-- 0x0d09
		"11111110",	-- 0x0d0a
		"11011010",	-- 0x0d0b
		"01001110",	-- 0x0d0c
		"10110010",	-- 0x0d0d
		"00000001",	-- 0x0d0e
		"11010101",	-- 0x0d0f
		"00110101",	-- 0x0d10
		"00011001",	-- 0x0d11
		"00000010",	-- 0x0d12
		"01110010",	-- 0x0d13
		"10111010",	-- 0x0d14
		"00110111",	-- 0x0d15
		"00010110",	-- 0x0d16
		"00011001",	-- 0x0d17
		"00110101",	-- 0x0d18
		"00110000",	-- 0x0d19
		"00010110",	-- 0x0d1a
		"01111001",	-- 0x0d1b
		"11000100",	-- 0x0d1c
		"01010111",	-- 0x0d1d
		"01000100",	-- 0x0d1e
		"00010011",	-- 0x0d1f
		"01111001",	-- 0x0d20
		"01000110",	-- 0x0d21
		"01010110",	-- 0x0d22
		"01000101",	-- 0x0d23
		"00001110",	-- 0x0d24
		"01111001",	-- 0x0d25
		"00001100",	-- 0x0d26
		"10111010",	-- 0x0d27
		"01000101",	-- 0x0d28
		"00001001",	-- 0x0d29
		"10110110",	-- 0x0d2a
		"00000001",	-- 0x0d2b
		"00001010",	-- 0x0d2c
		"00000100",	-- 0x0d2d
		"00000001",	-- 0x0d2e
		"11110011",	-- 0x0d2f
		"11010010",	-- 0x0d30
		"01110111",	-- 0x0d31
		"00110000",	-- 0x0d32
		"01000000",	-- 0x0d33
		"00110001",	-- 0x0d34
		"01110001",	-- 0x0d35
		"10010010",	-- 0x0d36
		"01000110",	-- 0x0d37
		"00101100",	-- 0x0d38
		"00110111",	-- 0x0d39
		"00010110",	-- 0x0d3a
		"00100111",	-- 0x0d3b
		"00110101",	-- 0x0d3c
		"00110000",	-- 0x0d3d
		"00100100",	-- 0x0d3e
		"01111001",	-- 0x0d3f
		"10110011",	-- 0x0d40
		"01010111",	-- 0x0d41
		"01000101",	-- 0x0d42
		"00100001",	-- 0x0d43
		"10010110",	-- 0x0d44
		"01010111",	-- 0x0d45
		"10001001",	-- 0x0d46
		"11110101",	-- 0x0d47
		"11000000",	-- 0x0d48
		"01000101",	-- 0x0d49
		"00000101",	-- 0x0d4a
		"01111001",	-- 0x0d4b
		"00111101",	-- 0x0d4c
		"10111010",	-- 0x0d4d
		"01000101",	-- 0x0d4e
		"00010101",	-- 0x0d4f
		"01111001",	-- 0x0d50
		"11100000",	-- 0x0d51
		"01010100",	-- 0x0d52
		"01000100",	-- 0x0d53
		"00010000",	-- 0x0d54
		"10000110",	-- 0x0d55
		"00000100",	-- 0x0d56
		"11100010",	-- 0x0d57
		"01111001",	-- 0x0d58
		"11011100",	-- 0x0d59
		"01010111",	-- 0x0d5a
		"01000100",	-- 0x0d5b
		"00000011",	-- 0x0d5c
		"10000110",	-- 0x0d5d
		"00001001",	-- 0x0d5e
		"11000100",	-- 0x0d5f
		"00000001",	-- 0x0d60
		"11110011",	-- 0x0d61
		"11010010",	-- 0x0d62
		"01110111",	-- 0x0d63
		"00110000",	-- 0x0d64
		"01100011",	-- 0x0d65
		"01000000",	-- 0x0d66
		"00100011",	-- 0x0d67
		"00110101",	-- 0x0d68
		"00010110",	-- 0x0d69
		"00011111",	-- 0x0d6a
		"00110111",	-- 0x0d6b
		"00010100",	-- 0x0d6c
		"00011100",	-- 0x0d6d
		"00110101",	-- 0x0d6e
		"01010110",	-- 0x0d6f
		"00011001",	-- 0x0d70
		"00110111",	-- 0x0d71
		"00010011",	-- 0x0d72
		"00001010",	-- 0x0d73
		"10001111",	-- 0x0d74
		"11000001",	-- 0x0d75
		"11010010",	-- 0x0d76
		"11011011",	-- 0x0d77
		"01011011",	-- 0x0d78
		"00000001",	-- 0x0d79
		"11000100",	-- 0x0d7a
		"01000100",	-- 0x0d7b
		"01000000",	-- 0x0d7c
		"00000110",	-- 0x0d7d
		"10001111",	-- 0x0d7e
		"11000001",	-- 0x0d7f
		"11011000",	-- 0x0d80
		"00000001",	-- 0x0d81
		"11000011",	-- 0x0d82
		"11101110",	-- 0x0d83
		"00000001",	-- 0x0d84
		"11000100",	-- 0x0d85
		"11001010",	-- 0x0d86
		"00000001",	-- 0x0d87
		"11110011",	-- 0x0d88
		"11010010",	-- 0x0d89
		"01100011",	-- 0x0d8a
		"01000000",	-- 0x0d8b
		"00101010",	-- 0x0d8c
		"11011010",	-- 0x0d8d
		"01011110",	-- 0x0d8e
		"01001010",	-- 0x0d8f
		"00000010",	-- 0x0d90
		"01110101",	-- 0x0d91
		"01110000",	-- 0x0d92
		"11001100",	-- 0x0d93
		"00001110",	-- 0x0d94
		"01001101",	-- 0x0d95
		"00011111",	-- 0x0d96
		"01111001",	-- 0x0d97
		"10100000",	-- 0x0d98
		"01011011",	-- 0x0d99
		"01000100",	-- 0x0d9a
		"00011010",	-- 0x0d9b
		"01111001",	-- 0x0d9c
		"00001110",	-- 0x0d9d
		"01010010",	-- 0x0d9e
		"01000101",	-- 0x0d9f
		"00010101",	-- 0x0da0
		"00110101",	-- 0x0da1
		"00010110",	-- 0x0da2
		"00010010",	-- 0x0da3
		"01110001",	-- 0x0da4
		"01110000",	-- 0x0da5
		"01000110",	-- 0x0da6
		"00001110",	-- 0x0da7
		"10001111",	-- 0x0da8
		"11000001",	-- 0x0da9
		"11111011",	-- 0x0daa
		"00000001",	-- 0x0dab
		"11000011",	-- 0x0dac
		"11101110",	-- 0x0dad
		"00000100",	-- 0x0dae
		"00000100",	-- 0x0daf
		"00000100",	-- 0x0db0
		"00000100",	-- 0x0db1
		"00000100",	-- 0x0db2
		"00000001",	-- 0x0db3
		"11110011",	-- 0x0db4
		"11010010",	-- 0x0db5
		"01100011",	-- 0x0db6
		"01000000",	-- 0x0db7
		"00010001",	-- 0x0db8
		"10000110",	-- 0x0db9
		"00000000",	-- 0x0dba
		"11111010",	-- 0x0dbb
		"01000000",	-- 0x0dbc
		"00001000",	-- 0x0dbd
		"01111001",	-- 0x0dbe
		"10001011",	-- 0x0dbf
		"01011100",	-- 0x0dc0
		"01000101",	-- 0x0dc1
		"00000110",	-- 0x0dc2
		"10000110",	-- 0x0dc3
		"00000000",	-- 0x0dc4
		"11111010",	-- 0x0dc5
		"00000001",	-- 0x0dc6
		"11110011",	-- 0x0dc7
		"11010010",	-- 0x0dc8
		"01100011",	-- 0x0dc9
		"11111010",	-- 0x0dca
		"00000001",	-- 0x0dcb
		"11010000",	-- 0x0dcc
		"10010010",	-- 0x0dcd
		"01001110",	-- 0x0dce
		"11001010",	-- 0x0dcf
		"10000000",	-- 0x0dd0
		"00110101",	-- 0x0dd1
		"01010100",	-- 0x0dd2
		"00000111",	-- 0x0dd3
		"01110101",	-- 0x0dd4
		"00011110",	-- 0x0dd5
		"10110010",	-- 0x0dd6
		"00000001",	-- 0x0dd7
		"00011100",	-- 0x0dd8
		"01000000",	-- 0x0dd9
		"00111111",	-- 0x0dda
		"01111001",	-- 0x0ddb
		"10001100",	-- 0x0ddc
		"01011001",	-- 0x0ddd
		"01000100",	-- 0x0dde
		"00110101",	-- 0x0ddf
		"01111001",	-- 0x0de0
		"00001010",	-- 0x0de1
		"01010010",	-- 0x0de2
		"01000101",	-- 0x0de3
		"00110000",	-- 0x0de4
		"00110111",	-- 0x0de5
		"01011101",	-- 0x0de6
		"00101101",	-- 0x0de7
		"01111001",	-- 0x0de8
		"11100100",	-- 0x0de9
		"01010111",	-- 0x0dea
		"01000011",	-- 0x0deb
		"00101011",	-- 0x0dec
		"01111001",	-- 0x0ded
		"01010000",	-- 0x0dee
		"01011001",	-- 0x0def
		"01000101",	-- 0x0df0
		"00100110",	-- 0x0df1
		"00110101",	-- 0x0df2
		"00011110",	-- 0x0df3
		"00100011",	-- 0x0df4
		"10001111",	-- 0x0df5
		"11000010",	-- 0x0df6
		"00000000",	-- 0x0df7
		"10010110",	-- 0x0df8
		"01010010",	-- 0x0df9
		"00000001",	-- 0x0dfa
		"11000011",	-- 0x0dfb
		"11110100",	-- 0x0dfc
		"11011100",	-- 0x0dfd
		"11010100",	-- 0x0dfe
		"01000100",	-- 0x0dff
		"00010111",	-- 0x0e00
		"11111010",	-- 0x0e01
		"00000010",	-- 0x0e02
		"00110111",	-- 0x0e03
		"11001100",	-- 0x0e04
		"00000100",	-- 0x0e05
		"01000101",	-- 0x0e06
		"00010000",	-- 0x0e07
		"01110101",	-- 0x0e08
		"00111110",	-- 0x0e09
		"10001111",	-- 0x0e0a
		"11000000",	-- 0x0e0b
		"11101110",	-- 0x0e0c
		"10000001",	-- 0x0e0d
		"00010100",	-- 0x0e0e
		"00111110",	-- 0x0e0f
		"10010110",	-- 0x0e10
		"01011001",	-- 0x0e11
		"00000001",	-- 0x0e12
		"11000100",	-- 0x0e13
		"10000110",	-- 0x0e14
		"10110010",	-- 0x0e15
		"00000001",	-- 0x0e16
		"00011100",	-- 0x0e17
		"01110111",	-- 0x0e18
		"00011110",	-- 0x0e19
		"11111010",	-- 0x0e1a
		"00000001",	-- 0x0e1b
		"00011100",	-- 0x0e1c
		"11001100",	-- 0x0e1d
		"10000000",	-- 0x0e1e
		"01000110",	-- 0x0e1f
		"00000110",	-- 0x0e20
		"01110001",	-- 0x0e21
		"00111110",	-- 0x0e22
		"01000110",	-- 0x0e23
		"00000010",	-- 0x0e24
		"01110010",	-- 0x0e25
		"11010100",	-- 0x0e26
		"01000000",	-- 0x0e27
		"01000011",	-- 0x0e28
		"11111010",	-- 0x0e29
		"00000001",	-- 0x0e2a
		"00011100",	-- 0x0e2b
		"01001011",	-- 0x0e2c
		"00001101",	-- 0x0e2d
		"11000000",	-- 0x0e2e
		"00010011",	-- 0x0e2f
		"11001100",	-- 0x0e30
		"10000000",	-- 0x0e31
		"01000101",	-- 0x0e32
		"00000100",	-- 0x0e33
		"11001010",	-- 0x0e34
		"10000000",	-- 0x0e35
		"01110010",	-- 0x0e36
		"11010100",	-- 0x0e37
		"10110010",	-- 0x0e38
		"00000001",	-- 0x0e39
		"00011100",	-- 0x0e3a
		"01100011",	-- 0x0e3b
		"11011010",	-- 0x0e3c
		"01011110",	-- 0x0e3d
		"11001100",	-- 0x0e3e
		"11110000",	-- 0x0e3f
		"01001101",	-- 0x0e40
		"00000111",	-- 0x0e41
		"11001100",	-- 0x0e42
		"11110100",	-- 0x0e43
		"01001101",	-- 0x0e44
		"00000101",	-- 0x0e45
		"01110101",	-- 0x0e46
		"01010100",	-- 0x0e47
		"10001100",	-- 0x0e48
		"01110111",	-- 0x0e49
		"01010100",	-- 0x0e4a
		"01011011",	-- 0x0e4b
		"11110100",	-- 0x0e4c
		"00000001",	-- 0x0e4d
		"00011101",	-- 0x0e4e
		"01001000",	-- 0x0e4f
		"00000111",	-- 0x0e50
		"01000101",	-- 0x0e51
		"00000011",	-- 0x0e52
		"11001010",	-- 0x0e53
		"10000000",	-- 0x0e54
		"10001100",	-- 0x0e55
		"11001010",	-- 0x0e56
		"01111111",	-- 0x0e57
		"10110010",	-- 0x0e58
		"00000001",	-- 0x0e59
		"00011110",	-- 0x0e5a
		"10110011",	-- 0x0e5b
		"00000001",	-- 0x0e5c
		"00011101",	-- 0x0e5d
		"11001100",	-- 0x0e5e
		"11110100",	-- 0x0e5f
		"01001101",	-- 0x0e60
		"00000111",	-- 0x0e61
		"11001100",	-- 0x0e62
		"11111000",	-- 0x0e63
		"01001101",	-- 0x0e64
		"00000101",	-- 0x0e65
		"01110101",	-- 0x0e66
		"01011101",	-- 0x0e67
		"10001100",	-- 0x0e68
		"01110111",	-- 0x0e69
		"01011101",	-- 0x0e6a
		"01100011",	-- 0x0e6b
		"01111001",	-- 0x0e6c
		"11011111",	-- 0x0e6d
		"01010111",	-- 0x0e6e
		"01000100",	-- 0x0e6f
		"00001000",	-- 0x0e70
		"01111001",	-- 0x0e71
		"11011010",	-- 0x0e72
		"01010111",	-- 0x0e73
		"01000100",	-- 0x0e74
		"00000101",	-- 0x0e75
		"01110101",	-- 0x0e76
		"01011110",	-- 0x0e77
		"10001100",	-- 0x0e78
		"01110111",	-- 0x0e79
		"01011110",	-- 0x0e7a
		"00110101",	-- 0x0e7b
		"01010110",	-- 0x0e7c
		"00000010",	-- 0x0e7d
		"01110010",	-- 0x0e7e
		"11010111",	-- 0x0e7f
		"01111001",	-- 0x0e80
		"00011111",	-- 0x0e81
		"11010111",	-- 0x0e82
		"01000100",	-- 0x0e83
		"00000101",	-- 0x0e84
		"01111001",	-- 0x0e85
		"01010010",	-- 0x0e86
		"01010010",	-- 0x0e87
		"01000101",	-- 0x0e88
		"00000010",	-- 0x0e89
		"01110101",	-- 0x0e8a
		"01111110",	-- 0x0e8b
		"01010011",	-- 0x0e8c
		"00110101",	-- 0x0e8d
		"00011001",	-- 0x0e8e
		"00111010",	-- 0x0e8f
		"00110101",	-- 0x0e90
		"00010110",	-- 0x0e91
		"00110111",	-- 0x0e92
		"00110111",	-- 0x0e93
		"01011110",	-- 0x0e94
		"00110100",	-- 0x0e95
		"00110101",	-- 0x0e96
		"01010110",	-- 0x0e97
		"00110001",	-- 0x0e98
		"01111001",	-- 0x0e99
		"00011001",	-- 0x0e9a
		"01011101",	-- 0x0e9b
		"01000101",	-- 0x0e9c
		"00101100",	-- 0x0e9d
		"11011010",	-- 0x0e9e
		"01000011",	-- 0x0e9f
		"11001110",	-- 0x0ea0
		"10011111",	-- 0x0ea1
		"01000110",	-- 0x0ea2
		"00100110",	-- 0x0ea3
		"01111001",	-- 0x0ea4
		"11111010",	-- 0x0ea5
		"01011101",	-- 0x0ea6
		"01000101",	-- 0x0ea7
		"00100100",	-- 0x0ea8
		"01111001",	-- 0x0ea9
		"00101100",	-- 0x0eaa
		"01011001",	-- 0x0eab
		"01000101",	-- 0x0eac
		"00011111",	-- 0x0ead
		"01111001",	-- 0x0eae
		"11110110",	-- 0x0eaf
		"01011110",	-- 0x0eb0
		"01001110",	-- 0x0eb1
		"00011010",	-- 0x0eb2
		"01111001",	-- 0x0eb3
		"01001000",	-- 0x0eb4
		"01010010",	-- 0x0eb5
		"01000010",	-- 0x0eb6
		"00010101",	-- 0x0eb7
		"11111010",	-- 0x0eb8
		"00000010",	-- 0x0eb9
		"00001000",	-- 0x0eba
		"11001100",	-- 0x0ebb
		"01100001",	-- 0x0ebc
		"01000011",	-- 0x0ebd
		"00001110",	-- 0x0ebe
		"01110001",	-- 0x0ebf
		"01111110",	-- 0x0ec0
		"01000110",	-- 0x0ec1
		"00001010",	-- 0x0ec2
		"10001111",	-- 0x0ec3
		"11000010",	-- 0x0ec4
		"00001001",	-- 0x0ec5
		"00000001",	-- 0x0ec6
		"11000011",	-- 0x0ec7
		"11110010",	-- 0x0ec8
		"01011011",	-- 0x0ec9
		"10110011",	-- 0x0eca
		"00000001",	-- 0x0ecb
		"00011111",	-- 0x0ecc
		"11011010",	-- 0x0ecd
		"01010010",	-- 0x0ece
		"10001111",	-- 0x0ecf
		"11000010",	-- 0x0ed0
		"00010100",	-- 0x0ed1
		"00000001",	-- 0x0ed2
		"11000011",	-- 0x0ed3
		"11110000",	-- 0x0ed4
		"10110001",	-- 0x0ed5
		"00000001",	-- 0x0ed6
		"00011111",	-- 0x0ed7
		"10110010",	-- 0x0ed8
		"00000001",	-- 0x0ed9
		"00100000",	-- 0x0eda
		"00000101",	-- 0x0edb
		"11111010",	-- 0x0edc
		"00000001",	-- 0x0edd
		"11011100",	-- 0x0ede
		"01011011",	-- 0x0edf
		"11000011",	-- 0x0ee0
		"11111101",	-- 0x0ee1
		"10110011",	-- 0x0ee2
		"00000001",	-- 0x0ee3
		"11011100",	-- 0x0ee4
		"00000111",	-- 0x0ee5
		"11001110",	-- 0x0ee6
		"00000010",	-- 0x0ee7
		"01000111",	-- 0x0ee8
		"00001011",	-- 0x0ee9
		"11111011",	-- 0x0eea
		"00000001",	-- 0x0eeb
		"00011111",	-- 0x0eec
		"11000101",	-- 0x0eed
		"00010011",	-- 0x0eee
		"01000100",	-- 0x0eef
		"00000001",	-- 0x0ef0
		"01010011",	-- 0x0ef1
		"10110011",	-- 0x0ef2
		"00000001",	-- 0x0ef3
		"00011111",	-- 0x0ef4
		"11111010",	-- 0x0ef5
		"00000001",	-- 0x0ef6
		"11011001",	-- 0x0ef7
		"10010010",	-- 0x0ef8
		"01001111",	-- 0x0ef9
		"11011010",	-- 0x0efa
		"01011111",	-- 0x0efb
		"01001011",	-- 0x0efc
		"00000010",	-- 0x0efd
		"01110010",	-- 0x0efe
		"10111011",	-- 0x0eff
		"00110101",	-- 0x0f00
		"00010110",	-- 0x0f01
		"00001110",	-- 0x0f02
		"00110101",	-- 0x0f03
		"10111100",	-- 0x0f04
		"00001011",	-- 0x0f05
		"00110101",	-- 0x0f06
		"11011100",	-- 0x0f07
		"00001000",	-- 0x0f08
		"01111001",	-- 0x0f09
		"00110001",	-- 0x0f0a
		"10111011",	-- 0x0f0b
		"01000101",	-- 0x0f0c
		"00000101",	-- 0x0f0d
		"01110111",	-- 0x0f0e
		"00011111",	-- 0x0f0f
		"10001100",	-- 0x0f10
		"01110101",	-- 0x0f11
		"00011111",	-- 0x0f12
		"01110101",	-- 0x0f13
		"10111111",	-- 0x0f14
		"11011010",	-- 0x0f15
		"01000011",	-- 0x0f16
		"11000010",	-- 0x0f17
		"10011111",	-- 0x0f18
		"01000111",	-- 0x0f19
		"00000011",	-- 0x0f1a
		"01110010",	-- 0x0f1b
		"11010010",	-- 0x0f1c
		"10001100",	-- 0x0f1d
		"01110010",	-- 0x0f1e
		"11010011",	-- 0x0f1f
		"00110101",	-- 0x0f20
		"11110110",	-- 0x0f21
		"00101110",	-- 0x0f22
		"00110101",	-- 0x0f23
		"00010110",	-- 0x0f24
		"00101011",	-- 0x0f25
		"11111010",	-- 0x0f26
		"00000010",	-- 0x0f27
		"01000010",	-- 0x0f28
		"11001110",	-- 0x0f29
		"01000000",	-- 0x0f2a
		"01000110",	-- 0x0f2b
		"00100100",	-- 0x0f2c
		"01111001",	-- 0x0f2d
		"00011111",	-- 0x0f2e
		"11010011",	-- 0x0f2f
		"01000100",	-- 0x0f30
		"00011111",	-- 0x0f31
		"01111001",	-- 0x0f32
		"11000100",	-- 0x0f33
		"01010111",	-- 0x0f34
		"01000101",	-- 0x0f35
		"00011010",	-- 0x0f36
		"10110110",	-- 0x0f37
		"00000001",	-- 0x0f38
		"00001010",	-- 0x0f39
		"10001001",	-- 0x0f3a
		"00000000",	-- 0x0f3b
		"10101111",	-- 0x0f3c
		"01000011",	-- 0x0f3d
		"00010010",	-- 0x0f3e
		"11011010",	-- 0x0f3f
		"01100000",	-- 0x0f40
		"01001010",	-- 0x0f41
		"00001110",	-- 0x0f42
		"00110101",	-- 0x0f43
		"11010011",	-- 0x0f44
		"00001011",	-- 0x0f45
		"00110101",	-- 0x0f46
		"01011000",	-- 0x0f47
		"00001000",	-- 0x0f48
		"00110101",	-- 0x0f49
		"01111101",	-- 0x0f4a
		"00000101",	-- 0x0f4b
		"01110111",	-- 0x0f4c
		"10111111",	-- 0x0f4d
		"00110101",	-- 0x0f4e
		"00011111",	-- 0x0f4f
		"00000101",	-- 0x0f50
		"01110101",	-- 0x0f51
		"00110110",	-- 0x0f52
		"00000011",	-- 0x0f53
		"11010000",	-- 0x0f54
		"01001111",	-- 0x0f55
		"01110111",	-- 0x0f56
		"00110110",	-- 0x0f57
		"00000101",	-- 0x0f58
		"11011010",	-- 0x0f59
		"01011111",	-- 0x0f5a
		"11011011",	-- 0x0f5b
		"01000100",	-- 0x0f5c
		"10011010",	-- 0x0f5d
		"01111000",	-- 0x0f5e
		"01110101",	-- 0x0f5f
		"10010100",	-- 0x0f60
		"00000111",	-- 0x0f61
		"00110111",	-- 0x0f62
		"01000000",	-- 0x0f63
		"00010011",	-- 0x0f64
		"01110101",	-- 0x0f65
		"10011111",	-- 0x0f66
		"10001111",	-- 0x0f67
		"11000010",	-- 0x0f68
		"00101101",	-- 0x0f69
		"01111001",	-- 0x0f6a
		"00011110",	-- 0x0f6b
		"01011101",	-- 0x0f6c
		"01000100",	-- 0x0f6d
		"00000101",	-- 0x0f6e
		"01111001",	-- 0x0f6f
		"00101111",	-- 0x0f70
		"01010000",	-- 0x0f71
		"01000101",	-- 0x0f72
		"00010100",	-- 0x0f73
		"00011101",	-- 0x0f74
		"00011101",	-- 0x0f75
		"01000000",	-- 0x0f76
		"00010000",	-- 0x0f77
		"10001111",	-- 0x0f78
		"11000010",	-- 0x0f79
		"00101001",	-- 0x0f7a
		"00110111",	-- 0x0f7b
		"01111111",	-- 0x0f7c
		"00001000",	-- 0x0f7d
		"00011101",	-- 0x0f7e
		"00011101",	-- 0x0f7f
		"00110111",	-- 0x0f80
		"10011111",	-- 0x0f81
		"00000011",	-- 0x0f82
		"10001111",	-- 0x0f83
		"00000001",	-- 0x0f84
		"00100001",	-- 0x0f85
		"01110111",	-- 0x0f86
		"10011111",	-- 0x0f87
		"00011011",	-- 0x0f88
		"10111010",	-- 0x0f89
		"00000001",	-- 0x0f8a
		"00100001",	-- 0x0f8b
		"10011110",	-- 0x0f8c
		"01111000",	-- 0x0f8d
		"01001010",	-- 0x0f8e
		"00000001",	-- 0x0f8f
		"01011010",	-- 0x0f90
		"10010010",	-- 0x0f91
		"01111010",	-- 0x0f92
		"10001111",	-- 0x0f93
		"11000010",	-- 0x0f94
		"00110001",	-- 0x0f95
		"01111001",	-- 0x0f96
		"00111001",	-- 0x0f97
		"01010000",	-- 0x0f98
		"01000101",	-- 0x0f99
		"00000011",	-- 0x0f9a
		"10001111",	-- 0x0f9b
		"11000010",	-- 0x0f9c
		"00111101",	-- 0x0f9d
		"00110101",	-- 0x0f9e
		"10011111",	-- 0x0f9f
		"00011001",	-- 0x0fa0
		"00011101",	-- 0x0fa1
		"00011101",	-- 0x0fa2
		"01101111",	-- 0x0fa3
		"11011011",	-- 0x0fa4
		"01011011",	-- 0x0fa5
		"00000001",	-- 0x0fa6
		"11000100",	-- 0x0fa7
		"01000100",	-- 0x0fa8
		"10110010",	-- 0x0fa9
		"00000001",	-- 0x0faa
		"00100011",	-- 0x0fab
		"11001010",	-- 0x0fac
		"00000101",	-- 0x0fad
		"01111111",	-- 0x0fae
		"00001101",	-- 0x0faf
		"11011011",	-- 0x0fb0
		"01011011",	-- 0x0fb1
		"00000001",	-- 0x0fb2
		"11000100",	-- 0x0fb3
		"01000100",	-- 0x0fb4
		"10110010",	-- 0x0fb5
		"00000001",	-- 0x0fb6
		"00100100",	-- 0x0fb7
		"01000000",	-- 0x0fb8
		"00000011",	-- 0x0fb9
		"00110111",	-- 0x0fba
		"01111111",	-- 0x0fbb
		"00000011",	-- 0x0fbc
		"10001111",	-- 0x0fbd
		"00000001",	-- 0x0fbe
		"00100011",	-- 0x0fbf
		"00011011",	-- 0x0fc0
		"10111010",	-- 0x0fc1
		"00000001",	-- 0x0fc2
		"00100011",	-- 0x0fc3
		"10011110",	-- 0x0fc4
		"01111000",	-- 0x0fc5
		"01001010",	-- 0x0fc6
		"00000001",	-- 0x0fc7
		"01011010",	-- 0x0fc8
		"10010010",	-- 0x0fc9
		"01111011",	-- 0x0fca
		"01110111",	-- 0x0fcb
		"01111111",	-- 0x0fcc
		"11001010",	-- 0x0fcd
		"00010000",	-- 0x0fce
		"11011110",	-- 0x0fcf
		"01111001",	-- 0x0fd0
		"01000111",	-- 0x0fd1
		"01001101",	-- 0x0fd2
		"00000001",	-- 0x0fd3
		"11011110",	-- 0x0fd4
		"01011010",	-- 0x0fd5
		"00000001",	-- 0x0fd6
		"11010001",	-- 0x0fd7
		"10000111",	-- 0x0fd8
		"11111010",	-- 0x0fd9
		"00000001",	-- 0x0fda
		"11010111",	-- 0x0fdb
		"11000110",	-- 0x0fdc
		"00000001",	-- 0x0fdd
		"10110010",	-- 0x0fde
		"00000001",	-- 0x0fdf
		"11010111",	-- 0x0fe0
		"01110010",	-- 0x0fe1
		"01111011",	-- 0x0fe2
		"00110111",	-- 0x0fe3
		"10011111",	-- 0x0fe4
		"01000000",	-- 0x0fe5
		"10001110",	-- 0x0fe6
		"11000010",	-- 0x0fe7
		"00101001",	-- 0x0fe8
		"10001111",	-- 0x0fe9
		"00000001",	-- 0x0fea
		"00100001",	-- 0x0feb
		"11001011",	-- 0x0fec
		"00000101",	-- 0x0fed
		"11011010",	-- 0x0fee
		"01111000",	-- 0x0fef
		"01001010",	-- 0x0ff0
		"00000100",	-- 0x0ff1
		"11001011",	-- 0x0ff2
		"00000101",	-- 0x0ff3
		"00011100",	-- 0x0ff4
		"00011101",	-- 0x0ff5
		"11101010",	-- 0x0ff6
		"10000000",	-- 0x0ff7
		"00001001",	-- 0x0ff8
		"01000101",	-- 0x0ff9
		"00000100",	-- 0x0ffa
		"11101100",	-- 0x0ffb
		"00000000",	-- 0x0ffc
		"01000100",	-- 0x0ffd
		"00000010",	-- 0x0ffe
		"11101010",	-- 0x0fff
		"00000000",	-- 0x1000
		"10000010",	-- 0x1001
		"10001111",	-- 0x1002
		"11000010",	-- 0x1003
		"00110001",	-- 0x1004
		"10001110",	-- 0x1005
		"00000001",	-- 0x1006
		"00100011",	-- 0x1007
		"11001011",	-- 0x1008
		"10100001",	-- 0x1009
		"11011010",	-- 0x100a
		"01111000",	-- 0x100b
		"01001010",	-- 0x100c
		"00000100",	-- 0x100d
		"11001011",	-- 0x100e
		"10100001",	-- 0x100f
		"00011100",	-- 0x1010
		"00011101",	-- 0x1011
		"11101010",	-- 0x1012
		"00000000",	-- 0x1013
		"00001001",	-- 0x1014
		"01000101",	-- 0x1015
		"00000100",	-- 0x1016
		"11101100",	-- 0x1017
		"10000000",	-- 0x1018
		"01000100",	-- 0x1019
		"00000001",	-- 0x101a
		"00011010",	-- 0x101b
		"10100010",	-- 0x101c
		"00000000",	-- 0x101d
		"01000000",	-- 0x101e
		"00000110",	-- 0x101f
		"01110010",	-- 0x1020
		"01111010",	-- 0x1021
		"01110001",	-- 0x1022
		"10110001",	-- 0x1023
		"01000110",	-- 0x1024
		"00100111",	-- 0x1025
		"10010110",	-- 0x1026
		"01100010",	-- 0x1027
		"10011110",	-- 0x1028
		"01111000",	-- 0x1029
		"01001010",	-- 0x102a
		"00001000",	-- 0x102b
		"10011000",	-- 0x102c
		"01111010",	-- 0x102d
		"01000100",	-- 0x102e
		"00001011",	-- 0x102f
		"01010010",	-- 0x1030
		"01010011",	-- 0x1031
		"01000000",	-- 0x1032
		"00000111",	-- 0x1033
		"10010111",	-- 0x1034
		"01111010",	-- 0x1035
		"01000100",	-- 0x1036
		"00000011",	-- 0x1037
		"10000110",	-- 0x1038
		"11111111",	-- 0x1039
		"11111111",	-- 0x103a
		"00110101",	-- 0x103b
		"00010011",	-- 0x103c
		"00000011",	-- 0x103d
		"00110111",	-- 0x103e
		"00110011",	-- 0x103f
		"00000101",	-- 0x1040
		"01111001",	-- 0x1041
		"00011111",	-- 0x1042
		"11010011",	-- 0x1043
		"01000101",	-- 0x1044
		"00011100",	-- 0x1045
		"10001111",	-- 0x1046
		"11000011",	-- 0x1047
		"10100001",	-- 0x1048
		"00100001",	-- 0x1049
		"10111111",	-- 0x104a
		"10011010",	-- 0x104b
		"01100010",	-- 0x104c
		"01000000",	-- 0x104d
		"00010101",	-- 0x104e
		"10000110",	-- 0x104f
		"10000000",	-- 0x1050
		"00000000",	-- 0x1051
		"10011010",	-- 0x1052
		"01100010",	-- 0x1053
		"01110101",	-- 0x1054
		"10010100",	-- 0x1055
		"01110111",	-- 0x1056
		"10110001",	-- 0x1057
		"11111010",	-- 0x1058
		"00000001",	-- 0x1059
		"11010111",	-- 0x105a
		"11000010",	-- 0x105b
		"11111110",	-- 0x105c
		"10110010",	-- 0x105d
		"00000001",	-- 0x105e
		"11010111",	-- 0x105f
		"01110101",	-- 0x1060
		"10011111",	-- 0x1061
		"01110101",	-- 0x1062
		"01111111",	-- 0x1063
		"10001111",	-- 0x1064
		"00000000",	-- 0x1065
		"10000101",	-- 0x1066
		"10001110",	-- 0x1067
		"11000011",	-- 0x1068
		"10100101",	-- 0x1069
		"00011011",	-- 0x106a
		"00011100",	-- 0x106b
		"00011100",	-- 0x106c
		"01101001",	-- 0x106d
		"00000001",	-- 0x106e
		"11000011",	-- 0x106f
		"11010111",	-- 0x1070
		"01101001",	-- 0x1071
		"01000101",	-- 0x1072
		"00000111",	-- 0x1073
		"10001101",	-- 0x1074
		"00000000",	-- 0x1075
		"10010101",	-- 0x1076
		"01000101",	-- 0x1077
		"11110001",	-- 0x1078
		"01000000",	-- 0x1079
		"00000011",	-- 0x107a
		"00000001",	-- 0x107b
		"11001000",	-- 0x107c
		"00001000",	-- 0x107d
		"01110101",	-- 0x107e
		"01011111",	-- 0x107f
		"00110111",	-- 0x1080
		"01010110",	-- 0x1081
		"00010010",	-- 0x1082
		"01111001",	-- 0x1083
		"00101000",	-- 0x1084
		"01011011",	-- 0x1085
		"01000100",	-- 0x1086
		"00100001",	-- 0x1087
		"01111001",	-- 0x1088
		"00010100",	-- 0x1089
		"01011011",	-- 0x108a
		"01000101",	-- 0x108b
		"00011100",	-- 0x108c
		"01111001",	-- 0x108d
		"00011000",	-- 0x108e
		"01010000",	-- 0x108f
		"01000101",	-- 0x1090
		"00010111",	-- 0x1091
		"01010010",	-- 0x1092
		"01000000",	-- 0x1093
		"00100101",	-- 0x1094
		"01111001",	-- 0x1095
		"10000000",	-- 0x1096
		"01011011",	-- 0x1097
		"01000100",	-- 0x1098
		"00001111",	-- 0x1099
		"01111001",	-- 0x109a
		"00011110",	-- 0x109b
		"01011011",	-- 0x109c
		"01000101",	-- 0x109d
		"00001010",	-- 0x109e
		"10010110",	-- 0x109f
		"01010000",	-- 0x10a0
		"11001100",	-- 0x10a1
		"01100001",	-- 0x10a2
		"01000100",	-- 0x10a3
		"00000100",	-- 0x10a4
		"11001100",	-- 0x10a5
		"00011000",	-- 0x10a6
		"01000100",	-- 0x10a7
		"00000110",	-- 0x10a8
		"00000011",	-- 0x10a9
		"11010001",	-- 0x10aa
		"01101101",	-- 0x10ab
		"00000011",	-- 0x10ac
		"00011111",	-- 0x10ad
		"00000110",	-- 0x10ae
		"10001111",	-- 0x10af
		"11010000",	-- 0x10b0
		"10101100",	-- 0x10b1
		"00000001",	-- 0x10b2
		"11000100",	-- 0x10b3
		"11001101",	-- 0x10b4
		"00000001",	-- 0x10b5
		"11000100",	-- 0x10b6
		"01110110",	-- 0x10b7
		"01010110",	-- 0x10b8
		"00010010",	-- 0x10b9
		"10001110",	-- 0x10ba
		"00000000",	-- 0x10bb
		"10000110",	-- 0x10bc
		"00001100",	-- 0x10bd
		"01111010",	-- 0x10be
		"01100111",	-- 0x10bf
		"11011100",	-- 0x10c0
		"01100111",	-- 0x10c1
		"01000111",	-- 0x10c2
		"00000010",	-- 0x10c3
		"01110010",	-- 0x10c4
		"01101001",	-- 0x10c5
		"00110101",	-- 0x10c6
		"00010000",	-- 0x10c7
		"11100000",	-- 0x10c8
		"00110111",	-- 0x10c9
		"00110110",	-- 0x10ca
		"11011101",	-- 0x10cb
		"01111001",	-- 0x10cc
		"11100011",	-- 0x10cd
		"01010111",	-- 0x10ce
		"01000011",	-- 0x10cf
		"11011000",	-- 0x10d0
		"00110101",	-- 0x10d1
		"01111011",	-- 0x10d2
		"11010101",	-- 0x10d3
		"11111010",	-- 0x10d4
		"00000010",	-- 0x10d5
		"00110001",	-- 0x10d6
		"11110110",	-- 0x10d7
		"00000010",	-- 0x10d8
		"00110010",	-- 0x10d9
		"11110110",	-- 0x10da
		"00000010",	-- 0x10db
		"00110011",	-- 0x10dc
		"11110110",	-- 0x10dd
		"00000010",	-- 0x10de
		"00110000",	-- 0x10df
		"11110110",	-- 0x10e0
		"00000010",	-- 0x10e1
		"00110110",	-- 0x10e2
		"01000110",	-- 0x10e3
		"11000100",	-- 0x10e4
		"01111001",	-- 0x10e5
		"10010011",	-- 0x10e6
		"01010110",	-- 0x10e7
		"01000101",	-- 0x10e8
		"10111111",	-- 0x10e9
		"00110101",	-- 0x10ea
		"10111001",	-- 0x10eb
		"10111100",	-- 0x10ec
		"11111010",	-- 0x10ed
		"00000001",	-- 0x10ee
		"11010001",	-- 0x10ef
		"11001110",	-- 0x10f0
		"00000100",	-- 0x10f1
		"01000110",	-- 0x10f2
		"10110101",	-- 0x10f3
		"11001110",	-- 0x10f4
		"00100000",	-- 0x10f5
		"01000111",	-- 0x10f6
		"00000100",	-- 0x10f7
		"11001110",	-- 0x10f8
		"00000001",	-- 0x10f9
		"01000111",	-- 0x10fa
		"10101101",	-- 0x10fb
		"01110111",	-- 0x10fc
		"01011111",	-- 0x10fd
		"00110111",	-- 0x10fe
		"00111111",	-- 0x10ff
		"01101000",	-- 0x1100
		"11001010",	-- 0x1101
		"00000110",	-- 0x1102
		"00110101",	-- 0x1103
		"01010110",	-- 0x1104
		"00000010",	-- 0x1105
		"11001010",	-- 0x1106
		"00000011",	-- 0x1107
		"11011100",	-- 0x1108
		"01101001",	-- 0x1109
		"01000010",	-- 0x110a
		"01011101",	-- 0x110b
		"11001011",	-- 0x110c
		"00000001",	-- 0x110d
		"01111001",	-- 0x110e
		"10001010",	-- 0x110f
		"01100100",	-- 0x1110
		"01000100",	-- 0x1111
		"00000110",	-- 0x1112
		"01010101",	-- 0x1113
		"01111001",	-- 0x1114
		"01110110",	-- 0x1115
		"01100100",	-- 0x1116
		"01000010",	-- 0x1117
		"01010000",	-- 0x1118
		"11100001",	-- 0x1119
		"00000000",	-- 0x111a
		"01101101",	-- 0x111b
		"00111100",	-- 0x111c
		"10000111",	-- 0x111d
		"11000011",	-- 0x111e
		"00100001",	-- 0x111f
		"00111111",	-- 0x1120
		"01111101",	-- 0x1121
		"00000001",	-- 0x1122
		"11000011",	-- 0x1123
		"11010111",	-- 0x1124
		"00000001",	-- 0x1125
		"11010001",	-- 0x1126
		"10011000",	-- 0x1127
		"01110101",	-- 0x1128
		"00011000",	-- 0x1129
		"11011011",	-- 0x112a
		"10000110",	-- 0x112b
		"11000101",	-- 0x112c
		"01011100",	-- 0x112d
		"01000100",	-- 0x112e
		"00000011",	-- 0x112f
		"01010101",	-- 0x1130
		"01110111",	-- 0x1131
		"00011000",	-- 0x1132
		"01010010",	-- 0x1133
		"10000101",	-- 0x1134
		"00000101",	-- 0x1135
		"10010011",	-- 0x1136
		"01111000",	-- 0x1137
		"01101001",	-- 0x1138
		"10001110",	-- 0x1139
		"00000000",	-- 0x113a
		"10010100",	-- 0x113b
		"00110011",	-- 0x113c
		"00000110",	-- 0x113d
		"01111001",	-- 0x113e
		"11011010",	-- 0x113f
		"01111001",	-- 0x1140
		"10010001",	-- 0x1141
		"01111000",	-- 0x1142
		"11010101",	-- 0x1143
		"01111000",	-- 0x1144
		"10000100",	-- 0x1145
		"00000000",	-- 0x1146
		"00110111",	-- 0x1147
		"00011000",	-- 0x1148
		"00000011",	-- 0x1149
		"00000001",	-- 0x114a
		"11000100",	-- 0x114b
		"11101100",	-- 0x114c
		"10000111",	-- 0x114d
		"00000000",	-- 0x114e
		"00100011",	-- 0x114f
		"10011010",	-- 0x1150
		"01111010",	-- 0x1151
		"11011011",	-- 0x1152
		"10000110",	-- 0x1153
		"01010010",	-- 0x1154
		"10011000",	-- 0x1155
		"01111010",	-- 0x1156
		"01001011",	-- 0x1157
		"00001001",	-- 0x1158
		"00000001",	-- 0x1159
		"11000100",	-- 0x115a
		"11100001",	-- 0x115b
		"11101101",	-- 0x115c
		"00000000",	-- 0x115d
		"01000011",	-- 0x115e
		"00000010",	-- 0x115f
		"01100001",	-- 0x1160
		"00110110",	-- 0x1161
		"00011110",	-- 0x1162
		"00011110",	-- 0x1163
		"01110000",	-- 0x1164
		"01111001",	-- 0x1165
		"01001010",	-- 0x1166
		"11010111",	-- 0x1167
		"01101001",	-- 0x1168
		"11101010",	-- 0x1169
		"00000000",	-- 0x116a
		"01000000",	-- 0x116b
		"00000111",	-- 0x116c
		"00110011",	-- 0x116d
		"11111111",	-- 0x116e
		"01100111",	-- 0x116f
		"01110010",	-- 0x1170
		"01101001",	-- 0x1171
		"11001010",	-- 0x1172
		"10000000",	-- 0x1173
		"00110101",	-- 0x1174
		"00110110",	-- 0x1175
		"00001000",	-- 0x1176
		"11001010",	-- 0x1177
		"10000000",	-- 0x1178
		"10010010",	-- 0x1179
		"01100100",	-- 0x117a
		"10010010",	-- 0x117b
		"01100001",	-- 0x117c
		"11001010",	-- 0x117d
		"00000000",	-- 0x117e
		"10110010",	-- 0x117f
		"00000010",	-- 0x1180
		"00011010",	-- 0x1181
		"01110101",	-- 0x1182
		"00111111",	-- 0x1183
		"00000011",	-- 0x1184
		"11010001",	-- 0x1185
		"11011101",	-- 0x1186
		"10010110",	-- 0x1187
		"01100001",	-- 0x1188
		"10010011",	-- 0x1189
		"01100001",	-- 0x118a
		"00001000",	-- 0x118b
		"00010100",	-- 0x118c
		"10010010",	-- 0x118d
		"01100100",	-- 0x118e
		"01110111",	-- 0x118f
		"00111111",	-- 0x1190
		"10000110",	-- 0x1191
		"01101001",	-- 0x1192
		"00000010",	-- 0x1193
		"00000001",	-- 0x1194
		"11000100",	-- 0x1195
		"10111001",	-- 0x1196
		"01100011",	-- 0x1197
		"11101010",	-- 0x1198
		"00000000",	-- 0x1199
		"00001001",	-- 0x119a
		"11100000",	-- 0x119b
		"00000001",	-- 0x119c
		"00000010",	-- 0x119d
		"10101010",	-- 0x119e
		"00000000",	-- 0x119f
		"01100011",	-- 0x11a0
		"11001011",	-- 0x11a1
		"10000000",	-- 0x11a2
		"00110111",	-- 0x11a3
		"00010010",	-- 0x11a4
		"00110110",	-- 0x11a5
		"00110111",	-- 0x11a6
		"01010110",	-- 0x11a7
		"00000100",	-- 0x11a8
		"11011011",	-- 0x11a9
		"10000110",	-- 0x11aa
		"01000000",	-- 0x11ab
		"00101111",	-- 0x11ac
		"10001111",	-- 0x11ad
		"11010000",	-- 0x11ae
		"10101100",	-- 0x11af
		"10010110",	-- 0x11b0
		"01010000",	-- 0x11b1
		"10001000",	-- 0x11b2
		"00000100",	-- 0x11b3
		"00001001",	-- 0x11b4
		"01000100",	-- 0x11b5
		"00000010",	-- 0x11b6
		"01010010",	-- 0x11b7
		"01010011",	-- 0x11b8
		"00000001",	-- 0x11b9
		"11000100",	-- 0x11ba
		"11001101",	-- 0x11bb
		"10001001",	-- 0x11bc
		"00001000",	-- 0x11bd
		"00011111",	-- 0x11be
		"01000011",	-- 0x11bf
		"00000100",	-- 0x11c0
		"10000111",	-- 0x11c1
		"00001000",	-- 0x11c2
		"00011111",	-- 0x11c3
		"00000100",	-- 0x11c4
		"00000001",	-- 0x11c5
		"11000100",	-- 0x11c6
		"01110110",	-- 0x11c7
		"01101101",	-- 0x11c8
		"00010010",	-- 0x11c9
		"10001111",	-- 0x11ca
		"00000000",	-- 0x11cb
		"10001000",	-- 0x11cc
		"00001101",	-- 0x11cd
		"11101010",	-- 0x11ce
		"10000000",	-- 0x11cf
		"11101011",	-- 0x11d0
		"10000010",	-- 0x11d1
		"00111111",	-- 0x11d2
		"01111101",	-- 0x11d3
		"01101111",	-- 0x11d4
		"00101110",	-- 0x11d5
		"01101001",	-- 0x11d6
		"00000001",	-- 0x11d7
		"11000100",	-- 0x11d8
		"01011100",	-- 0x11d9
		"01111111",	-- 0x11da
		"01011011",	-- 0x11db
		"01100011",	-- 0x11dc
		"11011010",	-- 0x11dd
		"01001110",	-- 0x11de
		"10110010",	-- 0x11df
		"00000001",	-- 0x11e0
		"11010000",	-- 0x11e1
		"11011010",	-- 0x11e2
		"01001111",	-- 0x11e3
		"10110010",	-- 0x11e4
		"00000001",	-- 0x11e5
		"11011001",	-- 0x11e6
		"01110001",	-- 0x11e7
		"11010001",	-- 0x11e8
		"01000110",	-- 0x11e9
		"00010010",	-- 0x11ea
		"10000110",	-- 0x11eb
		"11001101",	-- 0x11ec
		"00010100",	-- 0x11ed
		"00000001",	-- 0x11ee
		"11000100",	-- 0x11ef
		"10111001",	-- 0x11f0
		"00000001",	-- 0x11f1
		"11001001",	-- 0x11f2
		"00011010",	-- 0x11f3
		"00000001",	-- 0x11f4
		"11001011",	-- 0x11f5
		"00000000",	-- 0x11f6
		"00000001",	-- 0x11f7
		"11101100",	-- 0x11f8
		"00000111",	-- 0x11f9
		"00000001",	-- 0x11fa
		"11011110",	-- 0x11fb
		"01110001",	-- 0x11fc
		"01111001",	-- 0x11fd
		"01111010",	-- 0x11fe
		"11001000",	-- 0x11ff
		"01000101",	-- 0x1200
		"00001010",	-- 0x1201
		"01110010",	-- 0x1202
		"11001000",	-- 0x1203
		"10000110",	-- 0x1204
		"11101010",	-- 0x1205
		"00000101",	-- 0x1206
		"00000001",	-- 0x1207
		"11000100",	-- 0x1208
		"10111001",	-- 0x1209
		"01110110",	-- 0x120a
		"11101111",	-- 0x120b
		"01110001",	-- 0x120c
		"01010001",	-- 0x120d
		"01000111",	-- 0x120e
		"00000011",	-- 0x120f
		"00000011",	-- 0x1210
		"11010010",	-- 0x1211
		"11010010",	-- 0x1212
		"11011010",	-- 0x1213
		"01000011",	-- 0x1214
		"11000010",	-- 0x1215
		"10011111",	-- 0x1216
		"01000110",	-- 0x1217
		"00001111",	-- 0x1218
		"10110110",	-- 0x1219
		"00000001",	-- 0x121a
		"00100111",	-- 0x121b
		"10001001",	-- 0x121c
		"11111111",	-- 0x121d
		"11100111",	-- 0x121e
		"01001101",	-- 0x121f
		"00000111",	-- 0x1220
		"11111010",	-- 0x1221
		"00000010",	-- 0x1222
		"01000010",	-- 0x1223
		"11001110",	-- 0x1224
		"01000000",	-- 0x1225
		"01000111",	-- 0x1226
		"00000010",	-- 0x1227
		"01110010",	-- 0x1228
		"11010101",	-- 0x1229
		"11011010",	-- 0x122a
		"01101011",	-- 0x122b
		"01000110",	-- 0x122c
		"00001110",	-- 0x122d
		"10000110",	-- 0x122e
		"00001111",	-- 0x122f
		"00001100",	-- 0x1230
		"01111001",	-- 0x1231
		"00011110",	-- 0x1232
		"01011011",	-- 0x1233
		"01000101",	-- 0x1234
		"00000001",	-- 0x1235
		"01011010",	-- 0x1236
		"11111100",	-- 0x1237
		"00000001",	-- 0x1238
		"01000111",	-- 0x1239
		"01001110",	-- 0x123a
		"00000010",	-- 0x123b
		"01110110",	-- 0x123c
		"01101011",	-- 0x123d
		"00110101",	-- 0x123e
		"00110110",	-- 0x123f
		"00000011",	-- 0x1240
		"00000011",	-- 0x1241
		"11010010",	-- 0x1242
		"10111100",	-- 0x1243
		"10010110",	-- 0x1244
		"01010111",	-- 0x1245
		"10001001",	-- 0x1246
		"11100100",	-- 0x1247
		"11000000",	-- 0x1248
		"01000101",	-- 0x1249
		"01110001",	-- 0x124a
		"10001001",	-- 0x124b
		"11101111",	-- 0x124c
		"10000000",	-- 0x124d
		"01000100",	-- 0x124e
		"01101100",	-- 0x124f
		"11111010",	-- 0x1250
		"00000010",	-- 0x1251
		"00110001",	-- 0x1252
		"11110110",	-- 0x1253
		"00000010",	-- 0x1254
		"00110110",	-- 0x1255
		"01000110",	-- 0x1256
		"01100100",	-- 0x1257
		"01111001",	-- 0x1258
		"10000000",	-- 0x1259
		"01011011",	-- 0x125a
		"01000100",	-- 0x125b
		"01011111",	-- 0x125c
		"00110101",	-- 0x125d
		"00111001",	-- 0x125e
		"01011100",	-- 0x125f
		"11111010",	-- 0x1260
		"00000001",	-- 0x1261
		"01000111",	-- 0x1262
		"11001100",	-- 0x1263
		"11111110",	-- 0x1264
		"01001101",	-- 0x1265
		"01010101",	-- 0x1266
		"01111001",	-- 0x1267
		"10010011",	-- 0x1268
		"01010110",	-- 0x1269
		"01000101",	-- 0x126a
		"01010000",	-- 0x126b
		"01111001",	-- 0x126c
		"00111101",	-- 0x126d
		"11010101",	-- 0x126e
		"01000101",	-- 0x126f
		"01001011",	-- 0x1270
		"00110101",	-- 0x1271
		"01011100",	-- 0x1272
		"01001000",	-- 0x1273
		"11111010",	-- 0x1274
		"00000001",	-- 0x1275
		"11010001",	-- 0x1276
		"11001110",	-- 0x1277
		"00000100",	-- 0x1278
		"01000110",	-- 0x1279
		"01000001",	-- 0x127a
		"11001110",	-- 0x127b
		"00100000",	-- 0x127c
		"01000111",	-- 0x127d
		"00000100",	-- 0x127e
		"11001110",	-- 0x127f
		"00000001",	-- 0x1280
		"01000111",	-- 0x1281
		"00111001",	-- 0x1282
		"01111001",	-- 0x1283
		"00000110",	-- 0x1284
		"01101011",	-- 0x1285
		"01000011",	-- 0x1286
		"01001010",	-- 0x1287
		"11001010",	-- 0x1288
		"00000001",	-- 0x1289
		"11011011",	-- 0x128a
		"01011111",	-- 0x128b
		"01001010",	-- 0x128c
		"00000001",	-- 0x128d
		"01010100",	-- 0x128e
		"11010000",	-- 0x128f
		"01101100",	-- 0x1290
		"10010010",	-- 0x1291
		"01101100",	-- 0x1292
		"01111001",	-- 0x1293
		"00010001",	-- 0x1294
		"01101011",	-- 0x1295
		"01000101",	-- 0x1296
		"00111010",	-- 0x1297
		"00110101",	-- 0x1298
		"10110011",	-- 0x1299
		"00100001",	-- 0x129a
		"10010110",	-- 0x129b
		"10010110",	-- 0x129c
		"00110101",	-- 0x129d
		"00010010",	-- 0x129e
		"00000011",	-- 0x129f
		"10000110",	-- 0x12a0
		"00000000",	-- 0x12a1
		"11111111",	-- 0x12a2
		"01111001",	-- 0x12a3
		"10000100",	-- 0x12a4
		"01101100",	-- 0x12a5
		"01000100",	-- 0x12a6
		"00001100",	-- 0x12a7
		"01111001",	-- 0x12a8
		"01111100",	-- 0x12a9
		"01101100",	-- 0x12aa
		"01000010",	-- 0x12ab
		"00001111",	-- 0x12ac
		"01011000",	-- 0x12ad
		"01000111",	-- 0x12ae
		"00001100",	-- 0x12af
		"01010000",	-- 0x12b0
		"01010111",	-- 0x12b1
		"01000000",	-- 0x12b2
		"00000110",	-- 0x12b3
		"11001100",	-- 0x12b4
		"10000000",	-- 0x12b5
		"01000111",	-- 0x12b6
		"00000100",	-- 0x12b7
		"01010110",	-- 0x12b8
		"01010001",	-- 0x12b9
		"10011010",	-- 0x12ba
		"10010110",	-- 0x12bb
		"10000110",	-- 0x12bc
		"00000000",	-- 0x12bd
		"10000000",	-- 0x12be
		"10011010",	-- 0x12bf
		"01101011",	-- 0x12c0
		"01110101",	-- 0x12c1
		"10110011",	-- 0x12c2
		"01000000",	-- 0x12c3
		"00001101",	-- 0x12c4
		"11011011",	-- 0x12c5
		"10010110",	-- 0x12c6
		"10001111",	-- 0x12c7
		"11000011",	-- 0x12c8
		"10110111",	-- 0x12c9
		"00100001",	-- 0x12ca
		"10100000",	-- 0x12cb
		"01000100",	-- 0x12cc
		"00000011",	-- 0x12cd
		"00000001",	-- 0x12ce
		"11001000",	-- 0x12cf
		"00001000",	-- 0x12d0
		"01100011",	-- 0x12d1
		"00000001",	-- 0x12d2
		"11101010",	-- 0x12d3
		"00100010",	-- 0x12d4
		"00000001",	-- 0x12d5
		"11101000",	-- 0x12d6
		"01100101",	-- 0x12d7
		"11111010",	-- 0x12d8
		"00000001",	-- 0x12d9
		"11010111",	-- 0x12da
		"10010010",	-- 0x12db
		"01001110",	-- 0x12dc
		"11111010",	-- 0x12dd
		"00000001",	-- 0x12de
		"11011000",	-- 0x12df
		"10010010",	-- 0x12e0
		"01001111",	-- 0x12e1
		"00110101",	-- 0x12e2
		"01111010",	-- 0x12e3
		"00000011",	-- 0x12e4
		"01110101",	-- 0x12e5
		"01011111",	-- 0x12e6
		"10001100",	-- 0x12e7
		"01110111",	-- 0x12e8
		"01011111",	-- 0x12e9
		"00110101",	-- 0x12ea
		"11111001",	-- 0x12eb
		"00000011",	-- 0x12ec
		"01110101",	-- 0x12ed
		"01111111",	-- 0x12ee
		"10001100",	-- 0x12ef
		"01110111",	-- 0x12f0
		"01111111",	-- 0x12f1
		"00110101",	-- 0x12f2
		"00011010",	-- 0x12f3
		"00000011",	-- 0x12f4
		"01110101",	-- 0x12f5
		"00111111",	-- 0x12f6
		"10001100",	-- 0x12f7
		"01110111",	-- 0x12f8
		"00111111",	-- 0x12f9
		"00110101",	-- 0x12fa
		"10111001",	-- 0x12fb
		"00000011",	-- 0x12fc
		"01110101",	-- 0x12fd
		"10111111",	-- 0x12fe
		"10001100",	-- 0x12ff
		"01110111",	-- 0x1300
		"10111111",	-- 0x1301
		"00110101",	-- 0x1302
		"00111010",	-- 0x1303
		"00000011",	-- 0x1304
		"01110101",	-- 0x1305
		"10011111",	-- 0x1306
		"10001100",	-- 0x1307
		"01110111",	-- 0x1308
		"10011111",	-- 0x1309
		"00110101",	-- 0x130a
		"00011001",	-- 0x130b
		"00000011",	-- 0x130c
		"01110101",	-- 0x130d
		"00011111",	-- 0x130e
		"10001100",	-- 0x130f
		"01110111",	-- 0x1310
		"00011111",	-- 0x1311
		"00110101",	-- 0x1312
		"00010011",	-- 0x1313
		"00000010",	-- 0x1314
		"01110010",	-- 0x1315
		"11011100",	-- 0x1316
		"11011011",	-- 0x1317
		"10011010",	-- 0x1318
		"10001111",	-- 0x1319
		"11000011",	-- 0x131a
		"11000101",	-- 0x131b
		"00100001",	-- 0x131c
		"10010010",	-- 0x131d
		"01000100",	-- 0x131e
		"00000011",	-- 0x131f
		"00000001",	-- 0x1320
		"11001000",	-- 0x1321
		"00001000",	-- 0x1322
		"00110101",	-- 0x1323
		"00010110",	-- 0x1324
		"00010111",	-- 0x1325
		"01111001",	-- 0x1326
		"11100100",	-- 0x1327
		"01010111",	-- 0x1328
		"01000011",	-- 0x1329
		"00010010",	-- 0x132a
		"01111001",	-- 0x132b
		"00000010",	-- 0x132c
		"01011101",	-- 0x132d
		"01000100",	-- 0x132e
		"00001101",	-- 0x132f
		"11111010",	-- 0x1330
		"00000001",	-- 0x1331
		"11010101",	-- 0x1332
		"11001110",	-- 0x1333
		"00001000",	-- 0x1334
		"01000110",	-- 0x1335
		"00000110",	-- 0x1336
		"00110101",	-- 0x1337
		"10111111",	-- 0x1338
		"00000011",	-- 0x1339
		"01110111",	-- 0x133a
		"01011110",	-- 0x133b
		"10001100",	-- 0x133c
		"01110101",	-- 0x133d
		"01011110",	-- 0x133e
		"00110111",	-- 0x133f
		"01010110",	-- 0x1340
		"00001001",	-- 0x1341
		"00110101",	-- 0x1342
		"00111110",	-- 0x1343
		"00000110",	-- 0x1344
		"00110101",	-- 0x1345
		"11111110",	-- 0x1346
		"00000011",	-- 0x1347
		"00110111",	-- 0x1348
		"00011111",	-- 0x1349
		"00000010",	-- 0x134a
		"01110010",	-- 0x134b
		"11011011",	-- 0x134c
		"00110111",	-- 0x134d
		"00010110",	-- 0x134e
		"00010001",	-- 0x134f
		"01110010",	-- 0x1350
		"11011101",	-- 0x1351
		"11011010",	-- 0x1352
		"10011010",	-- 0x1353
		"00110101",	-- 0x1354
		"00010010",	-- 0x1355
		"00000010",	-- 0x1356
		"11001010",	-- 0x1357
		"01100110",	-- 0x1358
		"10000001",	-- 0x1359
		"00010000",	-- 0x135a
		"10000111",	-- 0x135b
		"00000000",	-- 0x135c
		"10100100",	-- 0x135d
		"10111010",	-- 0x135e
		"00000001",	-- 0x135f
		"10011011",	-- 0x1360
		"00110101",	-- 0x1361
		"00010110",	-- 0x1362
		"00001010",	-- 0x1363
		"01111001",	-- 0x1364
		"00101000",	-- 0x1365
		"01011101",	-- 0x1366
		"01000100",	-- 0x1367
		"00000101",	-- 0x1368
		"01111001",	-- 0x1369
		"10100000",	-- 0x136a
		"01011011",	-- 0x136b
		"01000101",	-- 0x136c
		"00000110",	-- 0x136d
		"10000110",	-- 0x136e
		"00001000",	-- 0x136f
		"10100100",	-- 0x1370
		"10111010",	-- 0x1371
		"00000001",	-- 0x1372
		"10100001",	-- 0x1373
		"01000000",	-- 0x1374
		"00001010",	-- 0x1375
		"10001111",	-- 0x1376
		"11000011",	-- 0x1377
		"00100011",	-- 0x1378
		"00000001",	-- 0x1379
		"11000011",	-- 0x137a
		"11101110",	-- 0x137b
		"10110010",	-- 0x137c
		"00000001",	-- 0x137d
		"10010001",	-- 0x137e
		"01100011",	-- 0x137f
		"01110001",	-- 0x1380
		"00110100",	-- 0x1381
		"01000110",	-- 0x1382
		"00100001",	-- 0x1383
		"00000001",	-- 0x1384
		"11010100",	-- 0x1385
		"11001001",	-- 0x1386
		"01000000",	-- 0x1387
		"00011100",	-- 0x1388
		"00000101",	-- 0x1389
		"01110101",	-- 0x138a
		"00100111",	-- 0x138b
		"10110110",	-- 0x138c
		"00000001",	-- 0x138d
		"10011000",	-- 0x138e
		"01000111",	-- 0x138f
		"00001000",	-- 0x1390
		"01110111",	-- 0x1391
		"00100110",	-- 0x1392
		"10010111",	-- 0x1393
		"00000100",	-- 0x1394
		"10011010",	-- 0x1395
		"00001010",	-- 0x1396
		"01110111",	-- 0x1397
		"00100111",	-- 0x1398
		"01110101",	-- 0x1399
		"00100110",	-- 0x139a
		"00000111",	-- 0x139b
		"00110101",	-- 0x139c
		"00111000",	-- 0x139d
		"00000011",	-- 0x139e
		"01110111",	-- 0x139f
		"00001001",	-- 0x13a0
		"10001100",	-- 0x13a1
		"01110101",	-- 0x13a2
		"00001001",	-- 0x13a3
		"01100011",	-- 0x13a4
		"00110111",	-- 0x13a5
		"00010000",	-- 0x13a6
		"00000011",	-- 0x13a7
		"00000011",	-- 0x13a8
		"11010100",	-- 0x13a9
		"11000110",	-- 0x13aa
		"00110101",	-- 0x13ab
		"11111110",	-- 0x13ac
		"00000011",	-- 0x13ad
		"00110101",	-- 0x13ae
		"10111111",	-- 0x13af
		"00000010",	-- 0x13b0
		"01110010",	-- 0x13b1
		"11101001",	-- 0x13b2
		"01010010",	-- 0x13b3
		"01010011",	-- 0x13b4
		"01111001",	-- 0x13b5
		"00111101",	-- 0x13b6
		"11000111",	-- 0x13b7
		"01000101",	-- 0x13b8
		"00000011",	-- 0x13b9
		"00000011",	-- 0x13ba
		"11010100",	-- 0x13bb
		"01110101",	-- 0x13bc
		"00110111",	-- 0x13bd
		"11110110",	-- 0x13be
		"00000110",	-- 0x13bf
		"10000110",	-- 0x13c0
		"00000010",	-- 0x13c1
		"00000000",	-- 0x13c2
		"00000011",	-- 0x13c3
		"11010100",	-- 0x13c4
		"01110101",	-- 0x13c5
		"00110111",	-- 0x13c6
		"10111111",	-- 0x13c7
		"01000101",	-- 0x13c8
		"01111001",	-- 0x13c9
		"11010010",	-- 0x13ca
		"01010111",	-- 0x13cb
		"01000101",	-- 0x13cc
		"01000000",	-- 0x13cd
		"00110111",	-- 0x13ce
		"01010110",	-- 0x13cf
		"00111101",	-- 0x13d0
		"10000110",	-- 0x13d1
		"00000010",	-- 0x13d2
		"00000000",	-- 0x13d3
		"00110101",	-- 0x13d4
		"11010110",	-- 0x13d5
		"00011000",	-- 0x13d6
		"10000110",	-- 0x13d7
		"00000010",	-- 0x13d8
		"00000000",	-- 0x13d9
		"01111001",	-- 0x13da
		"00100110",	-- 0x13db
		"11101001",	-- 0x13dc
		"01000100",	-- 0x13dd
		"00000011",	-- 0x13de
		"00000011",	-- 0x13df
		"11010100",	-- 0x13e0
		"01110101",	-- 0x13e1
		"11011011",	-- 0x13e2
		"10011010",	-- 0x13e3
		"00110101",	-- 0x13e4
		"00010010",	-- 0x13e5
		"00000010",	-- 0x13e6
		"11001011",	-- 0x13e7
		"01100110",	-- 0x13e8
		"01010010",	-- 0x13e9
		"00000110",	-- 0x13ea
		"00000110",	-- 0x13eb
		"00000011",	-- 0x13ec
		"11010100",	-- 0x13ed
		"01110101",	-- 0x13ee
		"01111001",	-- 0x13ef
		"00010111",	-- 0x13f0
		"11101001",	-- 0x13f1
		"01000100",	-- 0x13f2
		"00000110",	-- 0x13f3
		"00000001",	-- 0x13f4
		"11010100",	-- 0x13f5
		"10001001",	-- 0x13f6
		"00000011",	-- 0x13f7
		"11010100",	-- 0x13f8
		"10000000",	-- 0x13f9
		"01111001",	-- 0x13fa
		"10011001",	-- 0x13fb
		"11101001",	-- 0x13fc
		"01000101",	-- 0x13fd
		"01110110",	-- 0x13fe
		"00000001",	-- 0x13ff
		"11010100",	-- 0x1400
		"10010101",	-- 0x1401
		"10001000",	-- 0x1402
		"00000010",	-- 0x1403
		"00000000",	-- 0x1404
		"01000101",	-- 0x1405
		"00000010",	-- 0x1406
		"01010010",	-- 0x1407
		"01010011",	-- 0x1408
		"00000001",	-- 0x1409
		"11000100",	-- 0x140a
		"11101100",	-- 0x140b
		"01000000",	-- 0x140c
		"01110010",	-- 0x140d
		"01111001",	-- 0x140e
		"00111101",	-- 0x140f
		"11010000",	-- 0x1410
		"01000101",	-- 0x1411
		"00100001",	-- 0x1412
		"00110101",	-- 0x1413
		"01010110",	-- 0x1414
		"00011110",	-- 0x1415
		"01111001",	-- 0x1416
		"11010010",	-- 0x1417
		"01010111",	-- 0x1418
		"01000101",	-- 0x1419
		"00011001",	-- 0x141a
		"10001110",	-- 0x141b
		"01100001",	-- 0x141c
		"01010000",	-- 0x141d
		"11111011",	-- 0x141e
		"00000001",	-- 0x141f
		"01000100",	-- 0x1420
		"00000001",	-- 0x1421
		"11000101",	-- 0x1422
		"01001111",	-- 0x1423
		"00110111",	-- 0x1424
		"11111111",	-- 0x1425
		"00000011",	-- 0x1426
		"10001000",	-- 0x1427
		"00001010",	-- 0x1428
		"00111110",	-- 0x1429
		"10011001",	-- 0x142a
		"01010000",	-- 0x142b
		"01000010",	-- 0x142c
		"00000110",	-- 0x142d
		"01110111",	-- 0x142e
		"11111111",	-- 0x142f
		"01010010",	-- 0x1430
		"01010011",	-- 0x1431
		"01000000",	-- 0x1432
		"01000001",	-- 0x1433
		"01110101",	-- 0x1434
		"11111111",	-- 0x1435
		"10000110",	-- 0x1436
		"00000011",	-- 0x1437
		"00000000",	-- 0x1438
		"01111001",	-- 0x1439
		"00011000",	-- 0x143a
		"10110110",	-- 0x143b
		"01000101",	-- 0x143c
		"00001000",	-- 0x143d
		"10000110",	-- 0x143e
		"00000011",	-- 0x143f
		"00000000",	-- 0x1440
		"01111001",	-- 0x1441
		"00011000",	-- 0x1442
		"10110111",	-- 0x1443
		"01000100",	-- 0x1444
		"00000101",	-- 0x1445
		"00110101",	-- 0x1446
		"11010110",	-- 0x1447
		"00110111",	-- 0x1448
		"01000000",	-- 0x1449
		"00101010",	-- 0x144a
		"01100001",	-- 0x144b
		"00111100",	-- 0x144c
		"01101000",	-- 0x144d
		"01100001",	-- 0x144e
		"01000101",	-- 0x144f
		"10111000",	-- 0x1450
		"00000001",	-- 0x1451
		"10011101",	-- 0x1452
		"01000101",	-- 0x1453
		"00000010",	-- 0x1454
		"01010010",	-- 0x1455
		"01010011",	-- 0x1456
		"00000001",	-- 0x1457
		"11000100",	-- 0x1458
		"11101100",	-- 0x1459
		"00101110",	-- 0x145a
		"00110111",	-- 0x145b
		"11010110",	-- 0x145c
		"00010001",	-- 0x145d
		"00110101",	-- 0x145e
		"00111000",	-- 0x145f
		"00001010",	-- 0x1460
		"10111111",	-- 0x1461
		"00000001",	-- 0x1462
		"10011101",	-- 0x1463
		"10001101",	-- 0x1464
		"00000010",	-- 0x1465
		"00000000",	-- 0x1466
		"01000010",	-- 0x1467
		"00010100",	-- 0x1468
		"01000000",	-- 0x1469
		"00000100",	-- 0x146a
		"10101001",	-- 0x146b
		"00000000",	-- 0x146c
		"01000100",	-- 0x146d
		"00001110",	-- 0x146e
		"10110110",	-- 0x146f
		"00000001",	-- 0x1470
		"10011101",	-- 0x1471
		"01100001",	-- 0x1472
		"00101101",	-- 0x1473
		"01111110",	-- 0x1474
		"00000101",	-- 0x1475
		"00110101",	-- 0x1476
		"11011111",	-- 0x1477
		"00001000",	-- 0x1478
		"01110101",	-- 0x1479
		"00111000",	-- 0x147a
		"01000000",	-- 0x147b
		"00000110",	-- 0x147c
		"01100001",	-- 0x147d
		"00100010",	-- 0x147e
		"01111110",	-- 0x147f
		"00000101",	-- 0x1480
		"01110111",	-- 0x1481
		"00111000",	-- 0x1482
		"10111010",	-- 0x1483
		"00000001",	-- 0x1484
		"10011000",	-- 0x1485
		"00000111",	-- 0x1486
		"01000000",	-- 0x1487
		"00111101",	-- 0x1488
		"11011011",	-- 0x1489
		"01010110",	-- 0x148a
		"10001111",	-- 0x148b
		"11000011",	-- 0x148c
		"10000101",	-- 0x148d
		"00000001",	-- 0x148e
		"11000100",	-- 0x148f
		"01000100",	-- 0x1490
		"00000001",	-- 0x1491
		"11000100",	-- 0x1492
		"11001010",	-- 0x1493
		"01100011",	-- 0x1494
		"11011011",	-- 0x1495
		"01010110",	-- 0x1496
		"10001111",	-- 0x1497
		"11000011",	-- 0x1498
		"10001011",	-- 0x1499
		"00000001",	-- 0x149a
		"11000100",	-- 0x149b
		"01000100",	-- 0x149c
		"00000001",	-- 0x149d
		"11000100",	-- 0x149e
		"11001010",	-- 0x149f
		"01100011",	-- 0x14a0
		"10101001",	-- 0x14a1
		"00000000",	-- 0x14a2
		"01000101",	-- 0x14a3
		"00010100",	-- 0x14a4
		"00111110",	-- 0x14a5
		"00000100",	-- 0x14a6
		"00000100",	-- 0x14a7
		"01011000",	-- 0x14a8
		"01000110",	-- 0x14a9
		"00000101",	-- 0x14aa
		"11111101",	-- 0x14ab
		"00000001",	-- 0x14ac
		"10010100",	-- 0x14ad
		"01000101",	-- 0x14ae
		"00000111",	-- 0x14af
		"11111011",	-- 0x14b0
		"00000001",	-- 0x14b1
		"10010100",	-- 0x14b2
		"01010010",	-- 0x14b3
		"00000110",	-- 0x14b4
		"00000110",	-- 0x14b5
		"01000001",	-- 0x14b6
		"00111100",	-- 0x14b7
		"10001100",	-- 0x14b8
		"10100110",	-- 0x14b9
		"00000000",	-- 0x14ba
		"01100011",	-- 0x14bb
		"10001111",	-- 0x14bc
		"11000011",	-- 0x14bd
		"01110110",	-- 0x14be
		"00000001",	-- 0x14bf
		"11000011",	-- 0x14c0
		"11101110",	-- 0x14c1
		"10110010",	-- 0x14c2
		"00000001",	-- 0x14c3
		"10010100",	-- 0x14c4
		"01100011",	-- 0x14c5
		"00000011",	-- 0x14c6
		"11011001",	-- 0x14c7
		"00110001",	-- 0x14c8
		"01111001",	-- 0x14c9
		"00111101",	-- 0x14ca
		"11010000",	-- 0x14cb
		"01000100",	-- 0x14cc
		"00011100",	-- 0x14cd
		"10001111",	-- 0x14ce
		"11000011",	-- 0x14cf
		"00111000",	-- 0x14d0
		"00000001",	-- 0x14d1
		"11000011",	-- 0x14d2
		"11101110",	-- 0x14d3
		"01101000",	-- 0x14d4
		"10001111",	-- 0x14d5
		"11000011",	-- 0x14d6
		"01000101",	-- 0x14d7
		"11011010",	-- 0x14d8
		"01010100",	-- 0x14d9
		"00000001",	-- 0x14da
		"11000011",	-- 0x14db
		"11110000",	-- 0x14dc
		"00101110",	-- 0x14dd
		"10101001",	-- 0x14de
		"00000000",	-- 0x14df
		"01000100",	-- 0x14e0
		"00000010",	-- 0x14e1
		"10100110",	-- 0x14e2
		"00000000",	-- 0x14e3
		"01111110",	-- 0x14e4
		"00000001",	-- 0x14e5
		"11000100",	-- 0x14e6
		"11001100",	-- 0x14e7
		"01000000",	-- 0x14e8
		"00001010",	-- 0x14e9
		"10110110",	-- 0x14ea
		"00000001",	-- 0x14eb
		"10001111",	-- 0x14ec
		"10001000",	-- 0x14ed
		"00000000",	-- 0x14ee
		"00000001",	-- 0x14ef
		"01000100",	-- 0x14f0
		"00000010",	-- 0x14f1
		"01010010",	-- 0x14f2
		"01010011",	-- 0x14f3
		"10111010",	-- 0x14f4
		"00000001",	-- 0x14f5
		"10001111",	-- 0x14f6
		"01111001",	-- 0x14f7
		"00001100",	-- 0x14f8
		"10110001",	-- 0x14f9
		"01000100",	-- 0x14fa
		"00100110",	-- 0x14fb
		"01111001",	-- 0x14fc
		"00000101",	-- 0x14fd
		"01011101",	-- 0x14fe
		"01000101",	-- 0x14ff
		"00100001",	-- 0x1500
		"01111001",	-- 0x1501
		"01010000",	-- 0x1502
		"01011011",	-- 0x1503
		"01000100",	-- 0x1504
		"00011100",	-- 0x1505
		"01111001",	-- 0x1506
		"10001010",	-- 0x1507
		"01011100",	-- 0x1508
		"01000101",	-- 0x1509
		"00010111",	-- 0x150a
		"01110111",	-- 0x150b
		"10011110",	-- 0x150c
		"01111001",	-- 0x150d
		"11011100",	-- 0x150e
		"01010111",	-- 0x150f
		"01000101",	-- 0x1510
		"00010010",	-- 0x1511
		"11011011",	-- 0x1512
		"01010000",	-- 0x1513
		"10001111",	-- 0x1514
		"11000011",	-- 0x1515
		"01001100",	-- 0x1516
		"00000001",	-- 0x1517
		"11000100",	-- 0x1518
		"01000111",	-- 0x1519
		"00000001",	-- 0x151a
		"11000100",	-- 0x151b
		"11001010",	-- 0x151c
		"10111010",	-- 0x151d
		"00000001",	-- 0x151e
		"10010010",	-- 0x151f
		"01000000",	-- 0x1520
		"00010100",	-- 0x1521
		"01110101",	-- 0x1522
		"10011110",	-- 0x1523
		"00110101",	-- 0x1524
		"10011110",	-- 0x1525
		"00001111",	-- 0x1526
		"10110110",	-- 0x1527
		"00000001",	-- 0x1528
		"10010010",	-- 0x1529
		"01000111",	-- 0x152a
		"00001010",	-- 0x152b
		"10001000",	-- 0x152c
		"00000000",	-- 0x152d
		"00001000",	-- 0x152e
		"01000100",	-- 0x152f
		"00000010",	-- 0x1530
		"01010010",	-- 0x1531
		"01010011",	-- 0x1532
		"10111010",	-- 0x1533
		"00000001",	-- 0x1534
		"10010010",	-- 0x1535
		"01111001",	-- 0x1536
		"00111101",	-- 0x1537
		"11010000",	-- 0x1538
		"01000100",	-- 0x1539
		"00000101",	-- 0x153a
		"10000110",	-- 0x153b
		"00000011",	-- 0x153c
		"00000000",	-- 0x153d
		"01000000",	-- 0x153e
		"00001010",	-- 0x153f
		"10110110",	-- 0x1540
		"00000001",	-- 0x1541
		"10101001",	-- 0x1542
		"10001000",	-- 0x1543
		"00000000",	-- 0x1544
		"00000100",	-- 0x1545
		"01000100",	-- 0x1546
		"00000010",	-- 0x1547
		"01010010",	-- 0x1548
		"01010011",	-- 0x1549
		"10111010",	-- 0x154a
		"00000001",	-- 0x154b
		"10101001",	-- 0x154c
		"01111001",	-- 0x154d
		"00001111",	-- 0x154e
		"11010000",	-- 0x154f
		"01000010",	-- 0x1550
		"00001100",	-- 0x1551
		"11111010",	-- 0x1552
		"00000010",	-- 0x1553
		"00110110",	-- 0x1554
		"11001100",	-- 0x1555
		"00001101",	-- 0x1556
		"01000101",	-- 0x1557
		"00000101",	-- 0x1558
		"10000110",	-- 0x1559
		"00000010",	-- 0x155a
		"00000000",	-- 0x155b
		"01000000",	-- 0x155c
		"00000111",	-- 0x155d
		"01111001",	-- 0x155e
		"00111100",	-- 0x155f
		"11101010",	-- 0x1560
		"01000101",	-- 0x1561
		"00000101",	-- 0x1562
		"01010010",	-- 0x1563
		"01010011",	-- 0x1564
		"10111010",	-- 0x1565
		"00000001",	-- 0x1566
		"10101011",	-- 0x1567
		"01010010",	-- 0x1568
		"01010011",	-- 0x1569
		"00110111",	-- 0x156a
		"11010110",	-- 0x156b
		"00101110",	-- 0x156c
		"10001110",	-- 0x156d
		"11000011",	-- 0x156e
		"01110010",	-- 0x156f
		"00110111",	-- 0x1570
		"00111111",	-- 0x1571
		"00000011",	-- 0x1572
		"10001110",	-- 0x1573
		"11000011",	-- 0x1574
		"01110100",	-- 0x1575
		"00000001",	-- 0x1576
		"11010110",	-- 0x1577
		"00001010",	-- 0x1578
		"10110110",	-- 0x1579
		"00000001",	-- 0x157a
		"10101101",	-- 0x157b
		"00110111",	-- 0x157c
		"10011111",	-- 0x157d
		"00000111",	-- 0x157e
		"10000111",	-- 0x157f
		"00000000",	-- 0x1580
		"00000010",	-- 0x1581
		"01000101",	-- 0x1582
		"00010001",	-- 0x1583
		"01000000",	-- 0x1584
		"00000111",	-- 0x1585
		"10001000",	-- 0x1586
		"00000000",	-- 0x1587
		"00000010",	-- 0x1588
		"01000100",	-- 0x1589
		"00000010",	-- 0x158a
		"01010010",	-- 0x158b
		"01010011",	-- 0x158c
		"00111111",	-- 0x158d
		"00000001",	-- 0x158e
		"11000100",	-- 0x158f
		"11011101",	-- 0x1590
		"11101101",	-- 0x1591
		"00000000",	-- 0x1592
		"01000101",	-- 0x1593
		"00000101",	-- 0x1594
		"11001010",	-- 0x1595
		"00010000",	-- 0x1596
		"10100001",	-- 0x1597
		"00000000",	-- 0x1598
		"01000001",	-- 0x1599
		"00111101",	-- 0x159a
		"10111010",	-- 0x159b
		"00000001",	-- 0x159c
		"10101101",	-- 0x159d
		"10001110",	-- 0x159e
		"11000011",	-- 0x159f
		"01101100",	-- 0x15a0
		"01100001",	-- 0x15a1
		"01100111",	-- 0x15a2
		"11101010",	-- 0x15a3
		"00000000",	-- 0x15a4
		"00110111",	-- 0x15a5
		"11010110",	-- 0x15a6
		"00100110",	-- 0x15a7
		"01110101",	-- 0x15a8
		"00011000",	-- 0x15a9
		"10001110",	-- 0x15aa
		"11000011",	-- 0x15ab
		"01101110",	-- 0x15ac
		"00110111",	-- 0x15ad
		"00111111",	-- 0x15ae
		"00000011",	-- 0x15af
		"10001110",	-- 0x15b0
		"11000011",	-- 0x15b1
		"01110000",	-- 0x15b2
		"01100001",	-- 0x15b3
		"01010101",	-- 0x15b4
		"11100100",	-- 0x15b5
		"00000000",	-- 0x15b6
		"01000101",	-- 0x15b7
		"00000011",	-- 0x15b8
		"01110111",	-- 0x15b9
		"00011000",	-- 0x15ba
		"01000001",	-- 0x15bb
		"01010100",	-- 0x15bc
		"10000001",	-- 0x15bd
		"00010000",	-- 0x15be
		"00000001",	-- 0x15bf
		"11000100",	-- 0x15c0
		"11101001",	-- 0x15c1
		"10110111",	-- 0x15c2
		"00000001",	-- 0x15c3
		"10101101",	-- 0x15c4
		"01001010",	-- 0x15c5
		"00000010",	-- 0x15c6
		"01010010",	-- 0x15c7
		"01010011",	-- 0x15c8
		"10111010",	-- 0x15c9
		"00000001",	-- 0x15ca
		"10100111",	-- 0x15cb
		"11101010",	-- 0x15cc
		"00000000",	-- 0x15cd
		"10000001",	-- 0x15ce
		"00010000",	-- 0x15cf
		"10110111",	-- 0x15d0
		"00000001",	-- 0x15d1
		"10101101",	-- 0x15d2
		"10110111",	-- 0x15d3
		"00000001",	-- 0x15d4
		"10101001",	-- 0x15d5
		"10110111",	-- 0x15d6
		"00000001",	-- 0x15d7
		"10101011",	-- 0x15d8
		"10011010",	-- 0x15d9
		"01111000",	-- 0x15da
		"10001111",	-- 0x15db
		"11000011",	-- 0x15dc
		"10010001",	-- 0x15dd
		"00110111",	-- 0x15de
		"11011010",	-- 0x15df
		"00000001",	-- 0x15e0
		"00011101",	-- 0x15e1
		"00110111",	-- 0x15e2
		"11111010",	-- 0x15e3
		"00000010",	-- 0x15e4
		"00011101",	-- 0x15e5
		"00011101",	-- 0x15e6
		"11101010",	-- 0x15e7
		"10000000",	-- 0x15e8
		"10000001",	-- 0x15e9
		"00010000",	-- 0x15ea
		"10010111",	-- 0x15eb
		"01111000",	-- 0x15ec
		"10011010",	-- 0x15ed
		"01111000",	-- 0x15ee
		"10111001",	-- 0x15ef
		"00000001",	-- 0x15f0
		"10010101",	-- 0x15f1
		"01000111",	-- 0x15f2
		"00000010",	-- 0x15f3
		"01110010",	-- 0x15f4
		"11011110",	-- 0x15f5
		"10111010",	-- 0x15f6
		"00000001",	-- 0x15f7
		"10010101",	-- 0x15f8
		"10010110",	-- 0x15f9
		"01011001",	-- 0x15fa
		"10111000",	-- 0x15fb
		"00000001",	-- 0x15fc
		"10010101",	-- 0x15fd
		"01000100",	-- 0x15fe
		"00000010",	-- 0x15ff
		"01010010",	-- 0x1600
		"01010011",	-- 0x1601
		"00000001",	-- 0x1602
		"11000100",	-- 0x1603
		"11011101",	-- 0x1604
		"10110011",	-- 0x1605
		"00000001",	-- 0x1606
		"10010111",	-- 0x1607
		"01000000",	-- 0x1608
		"00001000",	-- 0x1609
		"00110101",	-- 0x160a
		"01011111",	-- 0x160b
		"00000011",	-- 0x160c
		"00110111",	-- 0x160d
		"01111111",	-- 0x160e
		"00000001",	-- 0x160f
		"00011100",	-- 0x1610
		"01100011",	-- 0x1611
		"00110101",	-- 0x1612
		"11010110",	-- 0x1613
		"00100010",	-- 0x1614
		"00110111",	-- 0x1615
		"01011110",	-- 0x1616
		"00011111",	-- 0x1617
		"01111001",	-- 0x1618
		"01011100",	-- 0x1619
		"11011011",	-- 0x161a
		"01000101",	-- 0x161b
		"00011010",	-- 0x161c
		"10001111",	-- 0x161d
		"11000011",	-- 0x161e
		"01010111",	-- 0x161f
		"11111011",	-- 0x1620
		"00000001",	-- 0x1621
		"10010111",	-- 0x1622
		"00011101",	-- 0x1623
		"11101101",	-- 0x1624
		"10000000",	-- 0x1625
		"01000010",	-- 0x1626
		"11111011",	-- 0x1627
		"11101011",	-- 0x1628
		"10000101",	-- 0x1629
		"01010010",	-- 0x162a
		"10110111",	-- 0x162b
		"00000001",	-- 0x162c
		"10011011",	-- 0x162d
		"10001000",	-- 0x162e
		"00000000",	-- 0x162f
		"10000000",	-- 0x1630
		"01000100",	-- 0x1631
		"00011110",	-- 0x1632
		"01010010",	-- 0x1633
		"01010011",	-- 0x1634
		"01000000",	-- 0x1635
		"00011010",	-- 0x1636
		"01110010",	-- 0x1637
		"11011110",	-- 0x1638
		"01110010",	-- 0x1639
		"11011101",	-- 0x163a
		"00110101",	-- 0x163b
		"00010110",	-- 0x163c
		"00010001",	-- 0x163d
		"11011010",	-- 0x163e
		"10011010",	-- 0x163f
		"00110101",	-- 0x1640
		"00010010",	-- 0x1641
		"00000010",	-- 0x1642
		"11001010",	-- 0x1643
		"01100110",	-- 0x1644
		"10000001",	-- 0x1645
		"00010000",	-- 0x1646
		"10111001",	-- 0x1647
		"00000001",	-- 0x1648
		"10011011",	-- 0x1649
		"01000011",	-- 0x164a
		"00000011",	-- 0x164b
		"10111010",	-- 0x164c
		"00000001",	-- 0x164d
		"10011011",	-- 0x164e
		"01000000",	-- 0x164f
		"00101110",	-- 0x1650
		"10011010",	-- 0x1651
		"01111000",	-- 0x1652
		"11011010",	-- 0x1653
		"10011010",	-- 0x1654
		"00110101",	-- 0x1655
		"00010010",	-- 0x1656
		"00000010",	-- 0x1657
		"11001010",	-- 0x1658
		"01100110",	-- 0x1659
		"10000001",	-- 0x165a
		"00010000",	-- 0x165b
		"00110111",	-- 0x165c
		"01011111",	-- 0x165d
		"00001001",	-- 0x165e
		"10001000",	-- 0x165f
		"00000000",	-- 0x1660
		"00000000",	-- 0x1661
		"00111110",	-- 0x1662
		"10000111",	-- 0x1663
		"00000001",	-- 0x1664
		"01001000",	-- 0x1665
		"01000000",	-- 0x1666
		"00000111",	-- 0x1667
		"10001000",	-- 0x1668
		"00000000",	-- 0x1669
		"00110011",	-- 0x166a
		"00111110",	-- 0x166b
		"10000111",	-- 0x166c
		"00000001",	-- 0x166d
		"01111011",	-- 0x166e
		"10011001",	-- 0x166f
		"01111000",	-- 0x1670
		"01000011",	-- 0x1671
		"00001001",	-- 0x1672
		"01110010",	-- 0x1673
		"11011101",	-- 0x1674
		"00111100",	-- 0x1675
		"10011001",	-- 0x1676
		"01111000",	-- 0x1677
		"01000100",	-- 0x1678
		"00000010",	-- 0x1679
		"10010110",	-- 0x167a
		"01111000",	-- 0x167b
		"10111010",	-- 0x167c
		"00000001",	-- 0x167d
		"10011011",	-- 0x167e
		"00110111",	-- 0x167f
		"11010110",	-- 0x1680
		"00100011",	-- 0x1681
		"10001111",	-- 0x1682
		"11000011",	-- 0x1683
		"01010100",	-- 0x1684
		"00000001",	-- 0x1685
		"11000100",	-- 0x1686
		"00111100",	-- 0x1687
		"10010010",	-- 0x1688
		"01111000",	-- 0x1689
		"10001111",	-- 0x168a
		"11000011",	-- 0x168b
		"01010010",	-- 0x168c
		"01010010",	-- 0x168d
		"00001101",	-- 0x168e
		"10110110",	-- 0x168f
		"00000001",	-- 0x1690
		"10100111",	-- 0x1691
		"00000100",	-- 0x1692
		"00000100",	-- 0x1693
		"01011000",	-- 0x1694
		"01000110",	-- 0x1695
		"00000100",	-- 0x1696
		"00000001",	-- 0x1697
		"11000100",	-- 0x1698
		"01011100",	-- 0x1699
		"10001100",	-- 0x169a
		"11101010",	-- 0x169b
		"10000001",	-- 0x169c
		"11010100",	-- 0x169d
		"01111000",	-- 0x169e
		"01000100",	-- 0x169f
		"00000001",	-- 0x16a0
		"01010010",	-- 0x16a1
		"10110010",	-- 0x16a2
		"00000001",	-- 0x16a3
		"10100000",	-- 0x16a4
		"00110111",	-- 0x16a5
		"11010110",	-- 0x16a6
		"00011110",	-- 0x16a7
		"00110111",	-- 0x16a8
		"01011110",	-- 0x16a9
		"00011011",	-- 0x16aa
		"01111001",	-- 0x16ab
		"01011100",	-- 0x16ac
		"11011011",	-- 0x16ad
		"01000101",	-- 0x16ae
		"00010110",	-- 0x16af
		"10001111",	-- 0x16b0
		"11000011",	-- 0x16b1
		"01100001",	-- 0x16b2
		"11111011",	-- 0x16b3
		"00000001",	-- 0x16b4
		"10010111",	-- 0x16b5
		"00011101",	-- 0x16b6
		"11101101",	-- 0x16b7
		"10000000",	-- 0x16b8
		"01000010",	-- 0x16b9
		"11111011",	-- 0x16ba
		"11101011",	-- 0x16bb
		"10000101",	-- 0x16bc
		"01010010",	-- 0x16bd
		"10110111",	-- 0x16be
		"00000001",	-- 0x16bf
		"10100001",	-- 0x16c0
		"10001000",	-- 0x16c1
		"00000000",	-- 0x16c2
		"10000000",	-- 0x16c3
		"01000000",	-- 0x16c4
		"00000011",	-- 0x16c5
		"10110110",	-- 0x16c6
		"00000001",	-- 0x16c7
		"10100001",	-- 0x16c8
		"10001001",	-- 0x16c9
		"00001010",	-- 0x16ca
		"01100110",	-- 0x16cb
		"01000100",	-- 0x16cc
		"00100001",	-- 0x16cd
		"00111110",	-- 0x16ce
		"11111010",	-- 0x16cf
		"00000001",	-- 0x16d0
		"10100000",	-- 0x16d1
		"10000001",	-- 0x16d2
		"00010000",	-- 0x16d3
		"10001000",	-- 0x16d4
		"00001000",	-- 0x16d5
		"10100100",	-- 0x16d6
		"01000101",	-- 0x16d7
		"00000010",	-- 0x16d8
		"01010010",	-- 0x16d9
		"01010011",	-- 0x16da
		"00000001",	-- 0x16db
		"11000100",	-- 0x16dc
		"11101100",	-- 0x16dd
		"10001001",	-- 0x16de
		"00000100",	-- 0x16df
		"00000000",	-- 0x16e0
		"01000100",	-- 0x16e1
		"00000011",	-- 0x16e2
		"10000110",	-- 0x16e3
		"00000100",	-- 0x16e4
		"00000000",	-- 0x16e5
		"10011010",	-- 0x16e6
		"01111000",	-- 0x16e7
		"10011100",	-- 0x16e8
		"01111000",	-- 0x16e9
		"01000011",	-- 0x16ea
		"00000110",	-- 0x16eb
		"00111100",	-- 0x16ec
		"01000000",	-- 0x16ed
		"00000011",	-- 0x16ee
		"10000110",	-- 0x16ef
		"00001010",	-- 0x16f0
		"01100110",	-- 0x16f1
		"10111010",	-- 0x16f2
		"00000001",	-- 0x16f3
		"10100001",	-- 0x16f4
		"11111010",	-- 0x16f5
		"00000001",	-- 0x16f6
		"10011010",	-- 0x16f7
		"01010110",	-- 0x16f8
		"10110010",	-- 0x16f9
		"00000001",	-- 0x16fa
		"10011010",	-- 0x16fb
		"00110111",	-- 0x16fc
		"00010010",	-- 0x16fd
		"00010111",	-- 0x16fe
		"01111001",	-- 0x16ff
		"01100110",	-- 0x1700
		"10011010",	-- 0x1701
		"01000100",	-- 0x1702
		"00010010",	-- 0x1703
		"10110110",	-- 0x1704
		"00000001",	-- 0x1705
		"10010101",	-- 0x1706
		"10000111",	-- 0x1707
		"00000111",	-- 0x1708
		"00000000",	-- 0x1709
		"00110111",	-- 0x170a
		"11010010",	-- 0x170b
		"00000101",	-- 0x170c
		"10001000",	-- 0x170d
		"00000001",	-- 0x170e
		"00000000",	-- 0x170f
		"01000101",	-- 0x1710
		"00000100",	-- 0x1711
		"10011001",	-- 0x1712
		"01110100",	-- 0x1713
		"01000010",	-- 0x1714
		"00000010",	-- 0x1715
		"01110010",	-- 0x1716
		"11011101",	-- 0x1717
		"01111001",	-- 0x1718
		"01011100",	-- 0x1719
		"11011101",	-- 0x171a
		"01000101",	-- 0x171b
		"00010011",	-- 0x171c
		"11011010",	-- 0x171d
		"10011110",	-- 0x171e
		"11000110",	-- 0x171f
		"00000001",	-- 0x1720
		"10010010",	-- 0x1721
		"10011110",	-- 0x1722
		"11001011",	-- 0x1723
		"01100110",	-- 0x1724
		"10110011",	-- 0x1725
		"00000001",	-- 0x1726
		"10001110",	-- 0x1727
		"10001110",	-- 0x1728
		"00000000",	-- 0x1729
		"10011010",	-- 0x172a
		"00000001",	-- 0x172b
		"11010001",	-- 0x172c
		"10011000",	-- 0x172d
		"01110010",	-- 0x172e
		"11011101",	-- 0x172f
		"00110101",	-- 0x1730
		"11110110",	-- 0x1731
		"00011111",	-- 0x1732
		"01111001",	-- 0x1733
		"11101000",	-- 0x1734
		"01010111",	-- 0x1735
		"01000101",	-- 0x1736
		"00011010",	-- 0x1737
		"11111010",	-- 0x1738
		"00000010",	-- 0x1739
		"00110001",	-- 0x173a
		"11110110",	-- 0x173b
		"00000010",	-- 0x173c
		"00110110",	-- 0x173d
		"01000110",	-- 0x173e
		"00010010",	-- 0x173f
		"01111001",	-- 0x1740
		"10010011",	-- 0x1741
		"01010110",	-- 0x1742
		"01000101",	-- 0x1743
		"00001101",	-- 0x1744
		"00110101",	-- 0x1745
		"01011111",	-- 0x1746
		"00001010",	-- 0x1747
		"10110110",	-- 0x1748
		"00000001",	-- 0x1749
		"10101011",	-- 0x174a
		"01000110",	-- 0x174b
		"00000101",	-- 0x174c
		"10110110",	-- 0x174d
		"00000001",	-- 0x174e
		"10001111",	-- 0x174f
		"01000111",	-- 0x1750
		"00000010",	-- 0x1751
		"01110010",	-- 0x1752
		"11011110",	-- 0x1753
		"01111001",	-- 0x1754
		"01011100",	-- 0x1755
		"11011110",	-- 0x1756
		"01000101",	-- 0x1757
		"00101011",	-- 0x1758
		"10110110",	-- 0x1759
		"00000001",	-- 0x175a
		"10010101",	-- 0x175b
		"10000111",	-- 0x175c
		"00001000",	-- 0x175d
		"00000000",	-- 0x175e
		"10011000",	-- 0x175f
		"01110100",	-- 0x1760
		"01000100",	-- 0x1761
		"00000011",	-- 0x1762
		"00000001",	-- 0x1763
		"11000100",	-- 0x1764
		"11101100",	-- 0x1765
		"10001001",	-- 0x1766
		"00000000",	-- 0x1767
		"01100000",	-- 0x1768
		"01000010",	-- 0x1769
		"00011001",	-- 0x176a
		"11011010",	-- 0x176b
		"10011010",	-- 0x176c
		"00110101",	-- 0x176d
		"00010010",	-- 0x176e
		"00000010",	-- 0x176f
		"11001010",	-- 0x1770
		"01100110",	-- 0x1771
		"10000001",	-- 0x1772
		"00010000",	-- 0x1773
		"10000111",	-- 0x1774
		"00000000",	-- 0x1775
		"01111011",	-- 0x1776
		"10111001",	-- 0x1777
		"00000001",	-- 0x1778
		"10011011",	-- 0x1779
		"01000101",	-- 0x177a
		"00001000",	-- 0x177b
		"10001000",	-- 0x177c
		"00000000",	-- 0x177d
		"01001000",	-- 0x177e
		"10111001",	-- 0x177f
		"00000001",	-- 0x1780
		"10011011",	-- 0x1781
		"01000011",	-- 0x1782
		"00000010",	-- 0x1783
		"01110010",	-- 0x1784
		"11100010",	-- 0x1785
		"00110111",	-- 0x1786
		"10111111",	-- 0x1787
		"00001000",	-- 0x1788
		"11011010",	-- 0x1789
		"10011110",	-- 0x178a
		"11000110",	-- 0x178b
		"00000001",	-- 0x178c
		"10010010",	-- 0x178d
		"10011110",	-- 0x178e
		"01000000",	-- 0x178f
		"00001011",	-- 0x1790
		"01111001",	-- 0x1791
		"10011001",	-- 0x1792
		"11100010",	-- 0x1793
		"01000101",	-- 0x1794
		"00000110",	-- 0x1795
		"11011010",	-- 0x1796
		"10011110",	-- 0x1797
		"11000010",	-- 0x1798
		"11111110",	-- 0x1799
		"10010010",	-- 0x179a
		"10011110",	-- 0x179b
		"11011010",	-- 0x179c
		"10011110",	-- 0x179d
		"11011011",	-- 0x179e
		"10011010",	-- 0x179f
		"00110101",	-- 0x17a0
		"00010010",	-- 0x17a1
		"00000100",	-- 0x17a2
		"11000010",	-- 0x17a3
		"11111110",	-- 0x17a4
		"11001011",	-- 0x17a5
		"01100110",	-- 0x17a6
		"01111001",	-- 0x17a7
		"00010001",	-- 0x17a8
		"01011101",	-- 0x17a9
		"01000100",	-- 0x17aa
		"00010000",	-- 0x17ab
		"11001110",	-- 0x17ac
		"00000001",	-- 0x17ad
		"01000110",	-- 0x17ae
		"00001100",	-- 0x17af
		"11111011",	-- 0x17b0
		"00000001",	-- 0x17b1
		"10001110",	-- 0x17b2
		"10001111",	-- 0x17b3
		"11000011",	-- 0x17b4
		"11000101",	-- 0x17b5
		"00100001",	-- 0x17b6
		"10010010",	-- 0x17b7
		"01000100",	-- 0x17b8
		"00000101",	-- 0x17b9
		"11001011",	-- 0x17ba
		"01100110",	-- 0x17bb
		"10110011",	-- 0x17bc
		"00000001",	-- 0x17bd
		"10001110",	-- 0x17be
		"01111001",	-- 0x17bf
		"01011100",	-- 0x17c0
		"11011110",	-- 0x17c1
		"01000101",	-- 0x17c2
		"01010001",	-- 0x17c3
		"11111011",	-- 0x17c4
		"00000001",	-- 0x17c5
		"10011010",	-- 0x17c6
		"01000111",	-- 0x17c7
		"00001010",	-- 0x17c8
		"00010011",	-- 0x17c9
		"00010011",	-- 0x17ca
		"01000110",	-- 0x17cb
		"01001000",	-- 0x17cc
		"11011010",	-- 0x17cd
		"10011110",	-- 0x17ce
		"11001110",	-- 0x17cf
		"00000001",	-- 0x17d0
		"01000111",	-- 0x17d1
		"01000010",	-- 0x17d2
		"11011010",	-- 0x17d3
		"10011010",	-- 0x17d4
		"10000001",	-- 0x17d5
		"00010000",	-- 0x17d6
		"00111110",	-- 0x17d7
		"11111010",	-- 0x17d8
		"00000001",	-- 0x17d9
		"10010111",	-- 0x17da
		"11011011",	-- 0x17db
		"10011010",	-- 0x17dc
		"10111100",	-- 0x17dd
		"00000001",	-- 0x17de
		"10011011",	-- 0x17df
		"01000111",	-- 0x17e0
		"00010111",	-- 0x17e1
		"01000101",	-- 0x17e2
		"00001011",	-- 0x17e3
		"11001100",	-- 0x17e4
		"01111010",	-- 0x17e5
		"01000101",	-- 0x17e6
		"00010001",	-- 0x17e7
		"11000101",	-- 0x17e8
		"00000001",	-- 0x17e9
		"01000100",	-- 0x17ea
		"00001101",	-- 0x17eb
		"01010011",	-- 0x17ec
		"01000000",	-- 0x17ed
		"00001010",	-- 0x17ee
		"11001100",	-- 0x17ef
		"10000110",	-- 0x17f0
		"01000010",	-- 0x17f1
		"00000110",	-- 0x17f2
		"11000001",	-- 0x17f3
		"00000001",	-- 0x17f4
		"01000100",	-- 0x17f5
		"00000010",	-- 0x17f6
		"11001011",	-- 0x17f7
		"11111111",	-- 0x17f8
		"11111010",	-- 0x17f9
		"00000001",	-- 0x17fa
		"10001110",	-- 0x17fb
		"11000000",	-- 0x17fc
		"00001000",	-- 0x17fd
		"10010010",	-- 0x17fe
		"01111000",	-- 0x17ff
		"11000100",	-- 0x1800
		"00001011",	-- 0x1801
		"10010010",	-- 0x1802
		"01111001",	-- 0x1803
		"10001111",	-- 0x1804
		"00000000",	-- 0x1805
		"01111000",	-- 0x1806
		"00000001",	-- 0x1807
		"11000011",	-- 0x1808
		"11010111",	-- 0x1809
		"10001111",	-- 0x180a
		"11000011",	-- 0x180b
		"11000101",	-- 0x180c
		"00100001",	-- 0x180d
		"10010010",	-- 0x180e
		"10001110",	-- 0x180f
		"00000000",	-- 0x1810
		"10011010",	-- 0x1811
		"00000001",	-- 0x1812
		"11010001",	-- 0x1813
		"10011000",	-- 0x1814
		"10010110",	-- 0x1815
		"01011001",	-- 0x1816
		"10111000",	-- 0x1817
		"00000001",	-- 0x1818
		"10100101",	-- 0x1819
		"01000111",	-- 0x181a
		"00010001",	-- 0x181b
		"00010100",	-- 0x181c
		"00010101",	-- 0x181d
		"00000001",	-- 0x181e
		"11000100",	-- 0x181f
		"11010101",	-- 0x1820
		"10001001",	-- 0x1821
		"00000000",	-- 0x1822
		"00000000",	-- 0x1823
		"01000110",	-- 0x1824
		"00000001",	-- 0x1825
		"01010111",	-- 0x1826
		"10110111",	-- 0x1827
		"00000001",	-- 0x1828
		"10100101",	-- 0x1829
		"10111010",	-- 0x182a
		"00000001",	-- 0x182b
		"10100101",	-- 0x182c
		"10011110",	-- 0x182d
		"01011001",	-- 0x182e
		"01111001",	-- 0x182f
		"00000010",	-- 0x1830
		"01011101",	-- 0x1831
		"01000101",	-- 0x1832
		"00011011",	-- 0x1833
		"01111001",	-- 0x1834
		"00010100",	-- 0x1835
		"01011001",	-- 0x1836
		"01000100",	-- 0x1837
		"00010001",	-- 0x1838
		"01111001",	-- 0x1839
		"00001101",	-- 0x183a
		"01011001",	-- 0x183b
		"01000101",	-- 0x183c
		"00010001",	-- 0x183d
		"10110110",	-- 0x183e
		"00000001",	-- 0x183f
		"10100101",	-- 0x1840
		"10011000",	-- 0x1841
		"01011001",	-- 0x1842
		"01000101",	-- 0x1843
		"00000101",	-- 0x1844
		"10001001",	-- 0x1845
		"00000010",	-- 0x1846
		"00000000",	-- 0x1847
		"01000100",	-- 0x1848
		"00000101",	-- 0x1849
		"10000110",	-- 0x184a
		"00000100",	-- 0x184b
		"00000000",	-- 0x184c
		"01000000",	-- 0x184d
		"00010100",	-- 0x184e
		"00111100",	-- 0x184f
		"10000111",	-- 0x1850
		"00000001",	-- 0x1851
		"00000000",	-- 0x1852
		"10111000",	-- 0x1853
		"00000001",	-- 0x1854
		"10100011",	-- 0x1855
		"01000100",	-- 0x1856
		"00000010",	-- 0x1857
		"01010010",	-- 0x1858
		"01010011",	-- 0x1859
		"00000110",	-- 0x185a
		"01000101",	-- 0x185b
		"00000011",	-- 0x185c
		"00000110",	-- 0x185d
		"01000100",	-- 0x185e
		"00000011",	-- 0x185f
		"10000110",	-- 0x1860
		"11111111",	-- 0x1861
		"11111111",	-- 0x1862
		"00001010",	-- 0x1863
		"00000001",	-- 0x1864
		"10100011",	-- 0x1865
		"00111110",	-- 0x1866
		"11001010",	-- 0x1867
		"01010000",	-- 0x1868
		"01111001",	-- 0x1869
		"00111101",	-- 0x186a
		"11010000",	-- 0x186b
		"01000101",	-- 0x186c
		"00100011",	-- 0x186d
		"00110111",	-- 0x186e
		"01010110",	-- 0x186f
		"00100000",	-- 0x1870
		"10000110",	-- 0x1871
		"00001000",	-- 0x1872
		"00000000",	-- 0x1873
		"00110111",	-- 0x1874
		"01011110",	-- 0x1875
		"00001000",	-- 0x1876
		"00110111",	-- 0x1877
		"00011110",	-- 0x1878
		"00000101",	-- 0x1879
		"11111010",	-- 0x187a
		"00000001",	-- 0x187b
		"10010111",	-- 0x187c
		"10000001",	-- 0x187d
		"00010000",	-- 0x187e
		"10001111",	-- 0x187f
		"11000010",	-- 0x1880
		"11111110",	-- 0x1881
		"00000001",	-- 0x1882
		"11000100",	-- 0x1883
		"10001010",	-- 0x1884
		"00110111",	-- 0x1885
		"01011110",	-- 0x1886
		"00000011",	-- 0x1887
		"00110101",	-- 0x1888
		"00011110",	-- 0x1889
		"00000110",	-- 0x188a
		"11001100",	-- 0x188b
		"01010000",	-- 0x188c
		"01000100",	-- 0x188d
		"00000010",	-- 0x188e
		"11001010",	-- 0x188f
		"01010000",	-- 0x1890
		"10110010",	-- 0x1891
		"00000001",	-- 0x1892
		"10011111",	-- 0x1893
		"00110111",	-- 0x1894
		"11010110",	-- 0x1895
		"00011001",	-- 0x1896
		"11011011",	-- 0x1897
		"10011010",	-- 0x1898
		"00110101",	-- 0x1899
		"00010010",	-- 0x189a
		"00000010",	-- 0x189b
		"11001011",	-- 0x189c
		"01100110",	-- 0x189d
		"01010010",	-- 0x189e
		"11110001",	-- 0x189f
		"00000001",	-- 0x18a0
		"10100000",	-- 0x18a1
		"10000000",	-- 0x18a2
		"00000000",	-- 0x18a3
		"00000110",	-- 0x18a4
		"00000110",	-- 0x18a5
		"00000110",	-- 0x18a6
		"00000110",	-- 0x18a7
		"10110111",	-- 0x18a8
		"00000001",	-- 0x18a9
		"10100001",	-- 0x18aa
		"10001000",	-- 0x18ab
		"00001000",	-- 0x18ac
		"00000000",	-- 0x18ad
		"01000000",	-- 0x18ae
		"00000011",	-- 0x18af
		"10110110",	-- 0x18b0
		"00000001",	-- 0x18b1
		"10011011",	-- 0x18b2
		"10110111",	-- 0x18b3
		"00000001",	-- 0x18b4
		"10001111",	-- 0x18b5
		"00000100",	-- 0x18b6
		"10011010",	-- 0x18b7
		"01111000",	-- 0x18b8
		"01010010",	-- 0x18b9
		"01010011",	-- 0x18ba
		"00110101",	-- 0x18bb
		"10011111",	-- 0x18bc
		"00000110",	-- 0x18bd
		"00110101",	-- 0x18be
		"01011111",	-- 0x18bf
		"00000011",	-- 0x18c0
		"00110111",	-- 0x18c1
		"01111111",	-- 0x18c2
		"00010100",	-- 0x18c3
		"10001111",	-- 0x18c4
		"11000011",	-- 0x18c5
		"01001010",	-- 0x18c6
		"00110111",	-- 0x18c7
		"11010110",	-- 0x18c8
		"00000001",	-- 0x18c9
		"00011101",	-- 0x18ca
		"00110111",	-- 0x18cb
		"11010000",	-- 0x18cc
		"00000111",	-- 0x18cd
		"00011101",	-- 0x18ce
		"00011101",	-- 0x18cf
		"00110101",	-- 0x18d0
		"11010010",	-- 0x18d1
		"00000010",	-- 0x18d2
		"00011101",	-- 0x18d3
		"00011101",	-- 0x18d4
		"11101011",	-- 0x18d5
		"10000000",	-- 0x18d6
		"00000110",	-- 0x18d7
		"10010111",	-- 0x18d8
		"01111000",	-- 0x18d9
		"10011010",	-- 0x18da
		"01111000",	-- 0x18db
		"11111011",	-- 0x18dc
		"00000001",	-- 0x18dd
		"10010001",	-- 0x18de
		"01010010",	-- 0x18df
		"00000110",	-- 0x18e0
		"00000110",	-- 0x18e1
		"10110111",	-- 0x18e2
		"00000001",	-- 0x18e3
		"10010010",	-- 0x18e4
		"00000110",	-- 0x18e5
		"10010111",	-- 0x18e6
		"01111000",	-- 0x18e7
		"00111110",	-- 0x18e8
		"00111100",	-- 0x18e9
		"00000100",	-- 0x18ea
		"11110001",	-- 0x18eb
		"00000001",	-- 0x18ec
		"10011111",	-- 0x18ed
		"10000000",	-- 0x18ee
		"00000000",	-- 0x18ef
		"10001000",	-- 0x18f0
		"00000000",	-- 0x18f1
		"01010000",	-- 0x18f2
		"01111001",	-- 0x18f3
		"11100100",	-- 0x18f4
		"01010111",	-- 0x18f5
		"01000100",	-- 0x18f6
		"00001000",	-- 0x18f7
		"00110111",	-- 0x18f8
		"01111110",	-- 0x18f9
		"00001010",	-- 0x18fa
		"01111001",	-- 0x18fb
		"11011111",	-- 0x18fc
		"01010111",	-- 0x18fd
		"01000101",	-- 0x18fe
		"00000101",	-- 0x18ff
		"01111001",	-- 0x1900
		"00011111",	-- 0x1901
		"11011100",	-- 0x1902
		"01000100",	-- 0x1903
		"00000011",	-- 0x1904
		"00000011",	-- 0x1905
		"11011001",	-- 0x1906
		"00101001",	-- 0x1907
		"01110111",	-- 0x1908
		"01111110",	-- 0x1909
		"10011010",	-- 0x190a
		"01111000",	-- 0x190b
		"01111001",	-- 0x190c
		"01111000",	-- 0x190d
		"01011011",	-- 0x190e
		"01000100",	-- 0x190f
		"00001000",	-- 0x1910
		"01111001",	-- 0x1911
		"01110000",	-- 0x1912
		"01011011",	-- 0x1913
		"01000100",	-- 0x1914
		"00000101",	-- 0x1915
		"01110101",	-- 0x1916
		"11011111",	-- 0x1917
		"10001100",	-- 0x1918
		"01110111",	-- 0x1919
		"11011111",	-- 0x191a
		"11011011",	-- 0x191b
		"01011011",	-- 0x191c
		"10001111",	-- 0x191d
		"11000011",	-- 0x191e
		"00011101",	-- 0x191f
		"00000001",	-- 0x1920
		"11000100",	-- 0x1921
		"01000111",	-- 0x1922
		"01011011",	-- 0x1923
		"01010010",	-- 0x1924
		"10010111",	-- 0x1925
		"01111000",	-- 0x1926
		"01000000",	-- 0x1927
		"00000100",	-- 0x1928
		"01110101",	-- 0x1929
		"01111110",	-- 0x192a
		"01110101",	-- 0x192b
		"11011111",	-- 0x192c
		"10111010",	-- 0x192d
		"00000001",	-- 0x192e
		"10011101",	-- 0x192f
		"01100011",	-- 0x1930
		"01110101",	-- 0x1931
		"00111110",	-- 0x1932
		"01110101",	-- 0x1933
		"11111110",	-- 0x1934
		"11011010",	-- 0x1935
		"01001110",	-- 0x1936
		"10110010",	-- 0x1937
		"00000001",	-- 0x1938
		"11010111",	-- 0x1939
		"11011010",	-- 0x193a
		"01001111",	-- 0x193b
		"10110010",	-- 0x193c
		"00000001",	-- 0x193d
		"11011000",	-- 0x193e
		"11111010",	-- 0x193f
		"00000001",	-- 0x1940
		"11010001",	-- 0x1941
		"10010010",	-- 0x1942
		"01001110",	-- 0x1943
		"00110111",	-- 0x1944
		"11011110",	-- 0x1945
		"00001101",	-- 0x1946
		"00110101",	-- 0x1947
		"10111110",	-- 0x1948
		"00001010",	-- 0x1949
		"01111001",	-- 0x194a
		"10001010",	-- 0x194b
		"01100100",	-- 0x194c
		"01000010",	-- 0x194d
		"00000101",	-- 0x194e
		"01111001",	-- 0x194f
		"01110110",	-- 0x1950
		"01100100",	-- 0x1951
		"01000100",	-- 0x1952
		"00000010",	-- 0x1953
		"01110010",	-- 0x1954
		"01101010",	-- 0x1955
		"01111001",	-- 0x1956
		"00011110",	-- 0x1957
		"11101010",	-- 0x1958
		"01000101",	-- 0x1959
		"00101011",	-- 0x195a
		"00110101",	-- 0x195b
		"10111001",	-- 0x195c
		"00101000",	-- 0x195d
		"11001010",	-- 0x195e
		"11100011",	-- 0x195f
		"00110111",	-- 0x1960
		"00111110",	-- 0x1961
		"00000010",	-- 0x1962
		"11001010",	-- 0x1963
		"11100001",	-- 0x1964
		"11011100",	-- 0x1965
		"01010111",	-- 0x1966
		"01000010",	-- 0x1967
		"00011101",	-- 0x1968
		"11111010",	-- 0x1969
		"00000010",	-- 0x196a
		"00110001",	-- 0x196b
		"11110110",	-- 0x196c
		"00000010",	-- 0x196d
		"00110000",	-- 0x196e
		"11110110",	-- 0x196f
		"00000010",	-- 0x1970
		"00110110",	-- 0x1971
		"01000110",	-- 0x1972
		"00010010",	-- 0x1973
		"00110101",	-- 0x1974
		"11110000",	-- 0x1975
		"00001111",	-- 0x1976
		"00110101",	-- 0x1977
		"00110110",	-- 0x1978
		"00010100",	-- 0x1979
		"11111010",	-- 0x197a
		"00000010",	-- 0x197b
		"01000010",	-- 0x197c
		"11001110",	-- 0x197d
		"01000000",	-- 0x197e
		"01000111",	-- 0x197f
		"00000101",	-- 0x1980
		"00000001",	-- 0x1981
		"11011011",	-- 0x1982
		"10010010",	-- 0x1983
		"01000000",	-- 0x1984
		"00000011",	-- 0x1985
		"00000001",	-- 0x1986
		"11011011",	-- 0x1987
		"10001100",	-- 0x1988
		"01110101",	-- 0x1989
		"00111110",	-- 0x198a
		"00000011",	-- 0x198b
		"11011100",	-- 0x198c
		"01110111",	-- 0x198d
		"01110111",	-- 0x198e
		"00111110",	-- 0x198f
		"01111001",	-- 0x1990
		"00011000",	-- 0x1991
		"10110100",	-- 0x1992
		"01000100",	-- 0x1993
		"00000011",	-- 0x1994
		"00000011",	-- 0x1995
		"11011010",	-- 0x1996
		"00010000",	-- 0x1997
		"01110010",	-- 0x1998
		"10110100",	-- 0x1999
		"10110110",	-- 0x199a
		"00000010",	-- 0x199b
		"00100110",	-- 0x199c
		"10011010",	-- 0x199d
		"01111000",	-- 0x199e
		"10110110",	-- 0x199f
		"00000010",	-- 0x19a0
		"00101000",	-- 0x19a1
		"10011010",	-- 0x19a2
		"01111010",	-- 0x19a3
		"10110110",	-- 0x19a4
		"00000001",	-- 0x19a5
		"10111110",	-- 0x19a6
		"00110111",	-- 0x19a7
		"00011110",	-- 0x19a8
		"00000110",	-- 0x19a9
		"00110111",	-- 0x19aa
		"01111110",	-- 0x19ab
		"00000011",	-- 0x19ac
		"10110110",	-- 0x19ad
		"00000001",	-- 0x19ae
		"11000000",	-- 0x19af
		"10001110",	-- 0x19b0
		"00011110",	-- 0x19b1
		"10111000",	-- 0x19b2
		"00000001",	-- 0x19b3
		"11000101",	-- 0x19b4
		"00000111",	-- 0x19b5
		"10111110",	-- 0x19b6
		"00000010",	-- 0x19b7
		"00101010",	-- 0x19b8
		"00000001",	-- 0x19b9
		"11000101",	-- 0x19ba
		"00000111",	-- 0x19bb
		"00111100",	-- 0x19bc
		"10011000",	-- 0x19bd
		"01111010",	-- 0x19be
		"01000011",	-- 0x19bf
		"00100010",	-- 0x19c0
		"00111110",	-- 0x19c1
		"11001010",	-- 0x19c2
		"11001000",	-- 0x19c3
		"00000001",	-- 0x19c4
		"11000101",	-- 0x19c5
		"01011011",	-- 0x19c6
		"10010110",	-- 0x19c7
		"01111000",	-- 0x19c8
		"00000001",	-- 0x19c9
		"11000101",	-- 0x19ca
		"10011011",	-- 0x19cb
		"10001001",	-- 0x19cc
		"00000000",	-- 0x19cd
		"11001000",	-- 0x19ce
		"01000101",	-- 0x19cf
		"00001001",	-- 0x19d0
		"10010110",	-- 0x19d1
		"01111000",	-- 0x19d2
		"10010111",	-- 0x19d3
		"01111010",	-- 0x19d4
		"00111110",	-- 0x19d5
		"11001011",	-- 0x19d6
		"11001000",	-- 0x19d7
		"01000000",	-- 0x19d8
		"00001100",	-- 0x19d9
		"01101101",	-- 0x19da
		"00110101",	-- 0x19db
		"00011110",	-- 0x19dc
		"00011100",	-- 0x19dd
		"10110110",	-- 0x19de
		"00000001",	-- 0x19df
		"10111110",	-- 0x19e0
		"01000000",	-- 0x19e1
		"00010011",	-- 0x19e2
		"01010011",	-- 0x19e3
		"10011110",	-- 0x19e4
		"01111010",	-- 0x19e5
		"01101101",	-- 0x19e6
		"01101110",	-- 0x19e7
		"10110110",	-- 0x19e8
		"00000010",	-- 0x19e9
		"00101010",	-- 0x19ea
		"10001110",	-- 0x19eb
		"00011110",	-- 0x19ec
		"10111000",	-- 0x19ed
		"00000001",	-- 0x19ee
		"11000101",	-- 0x19ef
		"00000111",	-- 0x19f0
		"00111100",	-- 0x19f1
		"01111110",	-- 0x19f2
		"00000001",	-- 0x19f3
		"11000101",	-- 0x19f4
		"10011011",	-- 0x19f5
		"10111010",	-- 0x19f6
		"00000001",	-- 0x19f7
		"11000000",	-- 0x19f8
		"00111110",	-- 0x19f9
		"01111100",	-- 0x19fa
		"10110010",	-- 0x19fb
		"00000001",	-- 0x19fc
		"10111101",	-- 0x19fd
		"11001100",	-- 0x19fe
		"11001000",	-- 0x19ff
		"01000101",	-- 0x1a00
		"00001110",	-- 0x1a01
		"00110101",	-- 0x1a02
		"00011110",	-- 0x1a03
		"00001011",	-- 0x1a04
		"00001010",	-- 0x1a05
		"00000001",	-- 0x1a06
		"10111110",	-- 0x1a07
		"01110111",	-- 0x1a08
		"10011110",	-- 0x1a09
		"00000001",	-- 0x1a0a
		"11011011",	-- 0x1a0b
		"10100011",	-- 0x1a0c
		"10111010",	-- 0x1a0d
		"00000001",	-- 0x1a0e
		"11000100",	-- 0x1a0f
		"01111001",	-- 0x1a10
		"01111010",	-- 0x1a11
		"10110101",	-- 0x1a12
		"01000100",	-- 0x1a13
		"00000010",	-- 0x1a14
		"01000000",	-- 0x1a15
		"01001001",	-- 0x1a16
		"01110010",	-- 0x1a17
		"10110101",	-- 0x1a18
		"00110101",	-- 0x1a19
		"00011110",	-- 0x1a1a
		"01000100",	-- 0x1a1b
		"00110111",	-- 0x1a1c
		"10111110",	-- 0x1a1d
		"01000001",	-- 0x1a1e
		"10110110",	-- 0x1a1f
		"00000001",	-- 0x1a20
		"10111110",	-- 0x1a21
		"10011110",	-- 0x1a22
		"01011111",	-- 0x1a23
		"01001011",	-- 0x1a24
		"00010011",	-- 0x1a25
		"01111001",	-- 0x1a26
		"01110110",	-- 0x1a27
		"01100010",	-- 0x1a28
		"01000011",	-- 0x1a29
		"00100010",	-- 0x1a2a
		"00111110",	-- 0x1a2b
		"11111010",	-- 0x1a2c
		"00000001",	-- 0x1a2d
		"10111101",	-- 0x1a2e
		"11001100",	-- 0x1a2f
		"11001000",	-- 0x1a30
		"01000100",	-- 0x1a31
		"00011011",	-- 0x1a32
		"00111100",	-- 0x1a33
		"10000111",	-- 0x1a34
		"00000000",	-- 0x1a35
		"00001100",	-- 0x1a36
		"01000000",	-- 0x1a37
		"00001100",	-- 0x1a38
		"01111001",	-- 0x1a39
		"01100110",	-- 0x1a3a
		"01100010",	-- 0x1a3b
		"01000100",	-- 0x1a3c
		"00001111",	-- 0x1a3d
		"10001000",	-- 0x1a3e
		"00000000",	-- 0x1a3f
		"00000010",	-- 0x1a40
		"01000100",	-- 0x1a41
		"00000010",	-- 0x1a42
		"01010010",	-- 0x1a43
		"01010011",	-- 0x1a44
		"10001111",	-- 0x1a45
		"11000011",	-- 0x1a46
		"11000001",	-- 0x1a47
		"00100001",	-- 0x1a48
		"10011111",	-- 0x1a49
		"10111010",	-- 0x1a4a
		"00000001",	-- 0x1a4b
		"10111110",	-- 0x1a4c
		"00111110",	-- 0x1a4d
		"11111010",	-- 0x1a4e
		"00000001",	-- 0x1a4f
		"10111101",	-- 0x1a50
		"11001100",	-- 0x1a51
		"11001000",	-- 0x1a52
		"01000100",	-- 0x1a53
		"00000011",	-- 0x1a54
		"00001010",	-- 0x1a55
		"00000001",	-- 0x1a56
		"11000000",	-- 0x1a57
		"10001100",	-- 0x1a58
		"00000000",	-- 0x1a59
		"01001101",	-- 0x1a5a
		"01000101",	-- 0x1a5b
		"00000011",	-- 0x1a5c
		"00000001",	-- 0x1a5d
		"11011100",	-- 0x1a5e
		"00111101",	-- 0x1a5f
		"00000011",	-- 0x1a60
		"11011100",	-- 0x1a61
		"01110111",	-- 0x1a62
		"01111001",	-- 0x1a63
		"00010100",	-- 0x1a64
		"01011001",	-- 0x1a65
		"01000100",	-- 0x1a66
		"00001000",	-- 0x1a67
		"01111001",	-- 0x1a68
		"00010110",	-- 0x1a69
		"01010000",	-- 0x1a6a
		"01000101",	-- 0x1a6b
		"00000011",	-- 0x1a6c
		"00110101",	-- 0x1a6d
		"01010110",	-- 0x1a6e
		"00000010",	-- 0x1a6f
		"01110010",	-- 0x1a70
		"11100100",	-- 0x1a71
		"00110111",	-- 0x1a72
		"01011110",	-- 0x1a73
		"00000111",	-- 0x1a74
		"01111001",	-- 0x1a75
		"01000000",	-- 0x1a76
		"11100100",	-- 0x1a77
		"01000101",	-- 0x1a78
		"00000010",	-- 0x1a79
		"01110101",	-- 0x1a7a
		"00011110",	-- 0x1a7b
		"00110101",	-- 0x1a7c
		"00011110",	-- 0x1a7d
		"01000000",	-- 0x1a7e
		"00110111",	-- 0x1a7f
		"00111110",	-- 0x1a80
		"00011111",	-- 0x1a81
		"01111001",	-- 0x1a82
		"00010100",	-- 0x1a83
		"01011001",	-- 0x1a84
		"01000100",	-- 0x1a85
		"00001101",	-- 0x1a86
		"01111001",	-- 0x1a87
		"00010110",	-- 0x1a88
		"01010000",	-- 0x1a89
		"01000101",	-- 0x1a8a
		"00001000",	-- 0x1a8b
		"00110111",	-- 0x1a8c
		"01010110",	-- 0x1a8d
		"00000101",	-- 0x1a8e
		"01110111",	-- 0x1a8f
		"11011110",	-- 0x1a90
		"00000011",	-- 0x1a91
		"11011011",	-- 0x1a92
		"00110100",	-- 0x1a93
		"10110110",	-- 0x1a94
		"00000001",	-- 0x1a95
		"10111110",	-- 0x1a96
		"10001001",	-- 0x1a97
		"00000000",	-- 0x1a98
		"10000000",	-- 0x1a99
		"01000100",	-- 0x1a9a
		"00010001",	-- 0x1a9b
		"00110101",	-- 0x1a9c
		"10111110",	-- 0x1a9d
		"00001001",	-- 0x1a9e
		"01000000",	-- 0x1a9f
		"00011001",	-- 0x1aa0
		"11111010",	-- 0x1aa1
		"00000010",	-- 0x1aa2
		"01000010",	-- 0x1aa3
		"11001110",	-- 0x1aa4
		"01000000",	-- 0x1aa5
		"01000110",	-- 0x1aa6
		"00010010",	-- 0x1aa7
		"00000001",	-- 0x1aa8
		"11011011",	-- 0x1aa9
		"01111001",	-- 0x1aaa
		"01000000",	-- 0x1aab
		"00001101",	-- 0x1aac
		"01110111",	-- 0x1aad
		"00011110",	-- 0x1aae
		"00000001",	-- 0x1aaf
		"11011100",	-- 0x1ab0
		"00111101",	-- 0x1ab1
		"10001001",	-- 0x1ab2
		"11000111",	-- 0x1ab3
		"10101110",	-- 0x1ab4
		"01000011",	-- 0x1ab5
		"00000011",	-- 0x1ab6
		"00000001",	-- 0x1ab7
		"11011011",	-- 0x1ab8
		"01110111",	-- 0x1ab9
		"01110101",	-- 0x1aba
		"11011110",	-- 0x1abb
		"00000011",	-- 0x1abc
		"11011011",	-- 0x1abd
		"01110100",	-- 0x1abe
		"01110101",	-- 0x1abf
		"11011110",	-- 0x1ac0
		"10110110",	-- 0x1ac1
		"00000001",	-- 0x1ac2
		"11000100",	-- 0x1ac3
		"01110101",	-- 0x1ac4
		"11111110",	-- 0x1ac5
		"01111001",	-- 0x1ac6
		"10110011",	-- 0x1ac7
		"01100100",	-- 0x1ac8
		"01000100",	-- 0x1ac9
		"00010000",	-- 0x1aca
		"01111001",	-- 0x1acb
		"01001101",	-- 0x1acc
		"01100100",	-- 0x1acd
		"01000010",	-- 0x1ace
		"11101010",	-- 0x1acf
		"01110111",	-- 0x1ad0
		"11111110",	-- 0x1ad1
		"10001000",	-- 0x1ad2
		"00000111",	-- 0x1ad3
		"10101110",	-- 0x1ad4
		"01000100",	-- 0x1ad5
		"00001100",	-- 0x1ad6
		"01010010",	-- 0x1ad7
		"01010011",	-- 0x1ad8
		"01000000",	-- 0x1ad9
		"00001000",	-- 0x1ada
		"10000111",	-- 0x1adb
		"00000111",	-- 0x1adc
		"10101110",	-- 0x1add
		"01000100",	-- 0x1ade
		"00000011",	-- 0x1adf
		"10000110",	-- 0x1ae0
		"11111111",	-- 0x1ae1
		"11111111",	-- 0x1ae2
		"10111010",	-- 0x1ae3
		"00000001",	-- 0x1ae4
		"11000100",	-- 0x1ae5
		"10010110",	-- 0x1ae6
		"01100010",	-- 0x1ae7
		"00110101",	-- 0x1ae8
		"11111110",	-- 0x1ae9
		"00011100",	-- 0x1aea
		"10001001",	-- 0x1aeb
		"00101001",	-- 0x1aec
		"01011100",	-- 0x1aed
		"01000100",	-- 0x1aee
		"00000101",	-- 0x1aef
		"10000110",	-- 0x1af0
		"00011010",	-- 0x1af1
		"00000000",	-- 0x1af2
		"01000000",	-- 0x1af3
		"00000011",	-- 0x1af4
		"10001000",	-- 0x1af5
		"00001111",	-- 0x1af6
		"01011100",	-- 0x1af7
		"10011010",	-- 0x1af8
		"01100010",	-- 0x1af9
		"11011010",	-- 0x1afa
		"01100100",	-- 0x1afb
		"11001100",	-- 0x1afc
		"00101001",	-- 0x1afd
		"01000100",	-- 0x1afe
		"00000011",	-- 0x1aff
		"11001010",	-- 0x1b00
		"00011010",	-- 0x1b01
		"10001100",	-- 0x1b02
		"11000100",	-- 0x1b03
		"00001111",	-- 0x1b04
		"01000000",	-- 0x1b05
		"00011010",	-- 0x1b06
		"10001001",	-- 0x1b07
		"11010110",	-- 0x1b08
		"10100100",	-- 0x1b09
		"01000101",	-- 0x1b0a
		"00000101",	-- 0x1b0b
		"10000110",	-- 0x1b0c
		"11100110",	-- 0x1b0d
		"00000000",	-- 0x1b0e
		"01000000",	-- 0x1b0f
		"00000011",	-- 0x1b10
		"10000111",	-- 0x1b11
		"00001111",	-- 0x1b12
		"01011100",	-- 0x1b13
		"10011010",	-- 0x1b14
		"01100010",	-- 0x1b15
		"11011010",	-- 0x1b16
		"01100100",	-- 0x1b17
		"11001100",	-- 0x1b18
		"11010111",	-- 0x1b19
		"01000101",	-- 0x1b1a
		"00000011",	-- 0x1b1b
		"11001010",	-- 0x1b1c
		"11100110",	-- 0x1b1d
		"10001100",	-- 0x1b1e
		"11000000",	-- 0x1b1f
		"00001111",	-- 0x1b20
		"10010010",	-- 0x1b21
		"01100100",	-- 0x1b22
		"00000001",	-- 0x1b23
		"11011100",	-- 0x1b24
		"00111101",	-- 0x1b25
		"00110101",	-- 0x1b26
		"11111110",	-- 0x1b27
		"00001000",	-- 0x1b28
		"10001001",	-- 0x1b29
		"11000111",	-- 0x1b2a
		"10101110",	-- 0x1b2b
		"01000011",	-- 0x1b2c
		"00000011",	-- 0x1b2d
		"00000001",	-- 0x1b2e
		"11011011",	-- 0x1b2f
		"01110111",	-- 0x1b30
		"00000011",	-- 0x1b31
		"11011011",	-- 0x1b32
		"01110100",	-- 0x1b33
		"00110101",	-- 0x1b34
		"10111110",	-- 0x1b35
		"00001010",	-- 0x1b36
		"00000001",	-- 0x1b37
		"11011011",	-- 0x1b38
		"01110101",	-- 0x1b39
		"01111001",	-- 0x1b3a
		"00000011",	-- 0x1b3b
		"01101010",	-- 0x1b3c
		"01000101",	-- 0x1b3d
		"00110101",	-- 0x1b3e
		"01110111",	-- 0x1b3f
		"10111110",	-- 0x1b40
		"10110110",	-- 0x1b41
		"00000001",	-- 0x1b42
		"11000100",	-- 0x1b43
		"10011110",	-- 0x1b44
		"01011111",	-- 0x1b45
		"01001011",	-- 0x1b46
		"00001111",	-- 0x1b47
		"01111001",	-- 0x1b48
		"10000101",	-- 0x1b49
		"01100010",	-- 0x1b4a
		"01000011",	-- 0x1b4b
		"00011001",	-- 0x1b4c
		"10000111",	-- 0x1b4d
		"00000000",	-- 0x1b4e
		"00010000",	-- 0x1b4f
		"01000100",	-- 0x1b50
		"00010100",	-- 0x1b51
		"10000110",	-- 0x1b52
		"11111111",	-- 0x1b53
		"11111111",	-- 0x1b54
		"01000000",	-- 0x1b55
		"00001111",	-- 0x1b56
		"01111001",	-- 0x1b57
		"01110110",	-- 0x1b58
		"01100010",	-- 0x1b59
		"01000100",	-- 0x1b5a
		"00001010",	-- 0x1b5b
		"00110101",	-- 0x1b5c
		"01111110",	-- 0x1b5d
		"00000111",	-- 0x1b5e
		"10001000",	-- 0x1b5f
		"00000000",	-- 0x1b60
		"00010000",	-- 0x1b61
		"01000100",	-- 0x1b62
		"00000010",	-- 0x1b63
		"01010010",	-- 0x1b64
		"01010011",	-- 0x1b65
		"10111010",	-- 0x1b66
		"00000001",	-- 0x1b67
		"11000100",	-- 0x1b68
		"10110110",	-- 0x1b69
		"00000001",	-- 0x1b6a
		"10111110",	-- 0x1b6b
		"10001001",	-- 0x1b6c
		"00000000",	-- 0x1b6d
		"01001101",	-- 0x1b6e
		"01000101",	-- 0x1b6f
		"00000011",	-- 0x1b70
		"00000001",	-- 0x1b71
		"11011100",	-- 0x1b72
		"00111101",	-- 0x1b73
		"01100011",	-- 0x1b74
		"01110101",	-- 0x1b75
		"01011110",	-- 0x1b76
		"01110101",	-- 0x1b77
		"00011110",	-- 0x1b78
		"10000110",	-- 0x1b79
		"11001100",	-- 0x1b7a
		"11001101",	-- 0x1b7b
		"10111010",	-- 0x1b7c
		"00000001",	-- 0x1b7d
		"11000010",	-- 0x1b7e
		"01110101",	-- 0x1b7f
		"10111110",	-- 0x1b80
		"01010010",	-- 0x1b81
		"01010011",	-- 0x1b82
		"10111010",	-- 0x1b83
		"00000001",	-- 0x1b84
		"10111110",	-- 0x1b85
		"10000110",	-- 0x1b86
		"11001100",	-- 0x1b87
		"11001101",	-- 0x1b88
		"10111010",	-- 0x1b89
		"00000001",	-- 0x1b8a
		"11000100",	-- 0x1b8b
		"01010010",	-- 0x1b8c
		"10110010",	-- 0x1b8d
		"00000001",	-- 0x1b8e
		"10111101",	-- 0x1b8f
		"01000000",	-- 0x1b90
		"00000101",	-- 0x1b91
		"11001010",	-- 0x1b92
		"11001000",	-- 0x1b93
		"10110010",	-- 0x1b94
		"00000001",	-- 0x1b95
		"10111101",	-- 0x1b96
		"01010010",	-- 0x1b97
		"01010011",	-- 0x1b98
		"10111010",	-- 0x1b99
		"00000001",	-- 0x1b9a
		"11000000",	-- 0x1b9b
		"10000110",	-- 0x1b9c
		"11001100",	-- 0x1b9d
		"11001101",	-- 0x1b9e
		"10111010",	-- 0x1b9f
		"00000001",	-- 0x1ba0
		"11000110",	-- 0x1ba1
		"01100011",	-- 0x1ba2
		"01110101",	-- 0x1ba3
		"00011000",	-- 0x1ba4
		"10111110",	-- 0x1ba5
		"00000001",	-- 0x1ba6
		"11000000",	-- 0x1ba7
		"00110101",	-- 0x1ba8
		"10011110",	-- 0x1ba9
		"00001010",	-- 0x1baa
		"10111100",	-- 0x1bab
		"00000001",	-- 0x1bac
		"10111110",	-- 0x1bad
		"01000110",	-- 0x1bae
		"00000101",	-- 0x1baf
		"10110110",	-- 0x1bb0
		"00000001",	-- 0x1bb1
		"11000100",	-- 0x1bb2
		"01000000",	-- 0x1bb3
		"00101001",	-- 0x1bb4
		"10110110",	-- 0x1bb5
		"00000001",	-- 0x1bb6
		"11000010",	-- 0x1bb7
		"10001000",	-- 0x1bb8
		"11001100",	-- 0x1bb9
		"11001101",	-- 0x1bba
		"01000100",	-- 0x1bbb
		"00000011",	-- 0x1bbc
		"00000001",	-- 0x1bbd
		"11000100",	-- 0x1bbe
		"11100111",	-- 0x1bbf
		"00000001",	-- 0x1bc0
		"11000101",	-- 0x1bc1
		"00000111",	-- 0x1bc2
		"00110101",	-- 0x1bc3
		"00011000",	-- 0x1bc4
		"00001010",	-- 0x1bc5
		"10000111",	-- 0x1bc6
		"11001100",	-- 0x1bc7
		"11001101",	-- 0x1bc8
		"01000100",	-- 0x1bc9
		"00010000",	-- 0x1bca
		"10000110",	-- 0x1bcb
		"11111111",	-- 0x1bcc
		"11111111",	-- 0x1bcd
		"01000000",	-- 0x1bce
		"00001011",	-- 0x1bcf
		"10001000",	-- 0x1bd0
		"11001100",	-- 0x1bd1
		"11001101",	-- 0x1bd2
		"01000101",	-- 0x1bd3
		"00000010",	-- 0x1bd4
		"01010010",	-- 0x1bd5
		"01010011",	-- 0x1bd6
		"01010100",	-- 0x1bd7
		"01010101",	-- 0x1bd8
		"10000100",	-- 0x1bd9
		"00000000",	-- 0x1bda
		"00110101",	-- 0x1bdb
		"10011110",	-- 0x1bdc
		"01011100",	-- 0x1bdd
		"10111001",	-- 0x1bde
		"00000001",	-- 0x1bdf
		"11001000",	-- 0x1be0
		"01000011",	-- 0x1be1
		"00001110",	-- 0x1be2
		"00110111",	-- 0x1be3
		"00011110",	-- 0x1be4
		"01001111",	-- 0x1be5
		"00110111",	-- 0x1be6
		"00111110",	-- 0x1be7
		"01001100",	-- 0x1be8
		"10111110",	-- 0x1be9
		"00000001",	-- 0x1bea
		"11000100",	-- 0x1beb
		"10111100",	-- 0x1bec
		"00000001",	-- 0x1bed
		"11001000",	-- 0x1bee
		"01000010",	-- 0x1bef
		"00110011",	-- 0x1bf0
		"01110111",	-- 0x1bf1
		"01111110",	-- 0x1bf2
		"10110110",	-- 0x1bf3
		"00000001",	-- 0x1bf4
		"11001000",	-- 0x1bf5
		"01101000",	-- 0x1bf6
		"10001000",	-- 0x1bf7
		"11001100",	-- 0x1bf8
		"11001101",	-- 0x1bf9
		"01010100",	-- 0x1bfa
		"01010101",	-- 0x1bfb
		"10000100",	-- 0x1bfc
		"00000000",	-- 0x1bfd
		"00111110",	-- 0x1bfe
		"10000110",	-- 0x1bff
		"11001100",	-- 0x1c00
		"11001101",	-- 0x1c01
		"10111000",	-- 0x1c02
		"00000001",	-- 0x1c03
		"11000010",	-- 0x1c04
		"01000010",	-- 0x1c05
		"00000101",	-- 0x1c06
		"10110110",	-- 0x1c07
		"00000001",	-- 0x1c08
		"10111110",	-- 0x1c09
		"01000000",	-- 0x1c0a
		"00001011",	-- 0x1c0b
		"00000001",	-- 0x1c0c
		"11000101",	-- 0x1c0d
		"10011011",	-- 0x1c0e
		"10001111",	-- 0x1c0f
		"11000011",	-- 0x1c10
		"11000001",	-- 0x1c11
		"00100001",	-- 0x1c12
		"10011111",	-- 0x1c13
		"10111010",	-- 0x1c14
		"00000001",	-- 0x1c15
		"11000000",	-- 0x1c16
		"01111110",	-- 0x1c17
		"00110101",	-- 0x1c18
		"00011110",	-- 0x1c19
		"00000110",	-- 0x1c1a
		"10111010",	-- 0x1c1b
		"00000001",	-- 0x1c1c
		"10111110",	-- 0x1c1d
		"00001010",	-- 0x1c1e
		"00000001",	-- 0x1c1f
		"11000100",	-- 0x1c20
		"00111100",	-- 0x1c21
		"01000000",	-- 0x1c22
		"00010011",	-- 0x1c23
		"00111110",	-- 0x1c24
		"11111010",	-- 0x1c25
		"00000001",	-- 0x1c26
		"10111101",	-- 0x1c27
		"01000111",	-- 0x1c28
		"00001010",	-- 0x1c29
		"11001100",	-- 0x1c2a
		"11001000",	-- 0x1c2b
		"01000100",	-- 0x1c2c
		"00000110",	-- 0x1c2d
		"10110110",	-- 0x1c2e
		"00000001",	-- 0x1c2f
		"10111110",	-- 0x1c30
		"10111010",	-- 0x1c31
		"00000001",	-- 0x1c32
		"11000000",	-- 0x1c33
		"00111100",	-- 0x1c34
		"01110101",	-- 0x1c35
		"01111110",	-- 0x1c36
		"10111010",	-- 0x1c37
		"00000001",	-- 0x1c38
		"11000110",	-- 0x1c39
		"01110101",	-- 0x1c3a
		"10011110",	-- 0x1c3b
		"01100011",	-- 0x1c3c
		"01110101",	-- 0x1c3d
		"00011000",	-- 0x1c3e
		"10110110",	-- 0x1c3f
		"00000001",	-- 0x1c40
		"11000100",	-- 0x1c41
		"10001000",	-- 0x1c42
		"11001100",	-- 0x1c43
		"11001101",	-- 0x1c44
		"01000100",	-- 0x1c45
		"00000011",	-- 0x1c46
		"00000001",	-- 0x1c47
		"11000100",	-- 0x1c48
		"11100111",	-- 0x1c49
		"00111110",	-- 0x1c4a
		"10110110",	-- 0x1c4b
		"00000001",	-- 0x1c4c
		"10111110",	-- 0x1c4d
		"00000001",	-- 0x1c4e
		"11000101",	-- 0x1c4f
		"10011011",	-- 0x1c50
		"00110101",	-- 0x1c51
		"00011000",	-- 0x1c52
		"00001010",	-- 0x1c53
		"10000111",	-- 0x1c54
		"11001100",	-- 0x1c55
		"11001101",	-- 0x1c56
		"01000100",	-- 0x1c57
		"00010000",	-- 0x1c58
		"10000110",	-- 0x1c59
		"11111111",	-- 0x1c5a
		"11111111",	-- 0x1c5b
		"01000000",	-- 0x1c5c
		"00001011",	-- 0x1c5d
		"10001000",	-- 0x1c5e
		"11001100",	-- 0x1c5f
		"11001101",	-- 0x1c60
		"01000101",	-- 0x1c61
		"00000010",	-- 0x1c62
		"01010010",	-- 0x1c63
		"01010011",	-- 0x1c64
		"01010100",	-- 0x1c65
		"01010101",	-- 0x1c66
		"10000100",	-- 0x1c67
		"00000000",	-- 0x1c68
		"10111010",	-- 0x1c69
		"00000001",	-- 0x1c6a
		"11000010",	-- 0x1c6b
		"10001001",	-- 0x1c6c
		"11000111",	-- 0x1c6d
		"10101110",	-- 0x1c6e
		"01000010",	-- 0x1c6f
		"00000011",	-- 0x1c70
		"01110111",	-- 0x1c71
		"01011110",	-- 0x1c72
		"10001100",	-- 0x1c73
		"01110101",	-- 0x1c74
		"01011110",	-- 0x1c75
		"01100011",	-- 0x1c76
		"11011010",	-- 0x1c77
		"01001110",	-- 0x1c78
		"10110010",	-- 0x1c79
		"00000001",	-- 0x1c7a
		"11010001",	-- 0x1c7b
		"11111010",	-- 0x1c7c
		"00000001",	-- 0x1c7d
		"11011010",	-- 0x1c7e
		"10010010",	-- 0x1c7f
		"01001111",	-- 0x1c80
		"01111001",	-- 0x1c81
		"00110100",	-- 0x1c82
		"01011001",	-- 0x1c83
		"01000100",	-- 0x1c84
		"00000010",	-- 0x1c85
		"01110101",	-- 0x1c86
		"00011111",	-- 0x1c87
		"01111001",	-- 0x1c88
		"00111100",	-- 0x1c89
		"01011001",	-- 0x1c8a
		"01000101",	-- 0x1c8b
		"00000010",	-- 0x1c8c
		"01110111",	-- 0x1c8d
		"00011111",	-- 0x1c8e
		"11011010",	-- 0x1c8f
		"11001001",	-- 0x1c90
		"00110101",	-- 0x1c91
		"10011001",	-- 0x1c92
		"00000011",	-- 0x1c93
		"00110101",	-- 0x1c94
		"01011010",	-- 0x1c95
		"00000111",	-- 0x1c96
		"11001100",	-- 0x1c97
		"00011000",	-- 0x1c98
		"01000100",	-- 0x1c99
		"00000011",	-- 0x1c9a
		"01010010",	-- 0x1c9b
		"10010010",	-- 0x1c9c
		"11001001",	-- 0x1c9d
		"00110111",	-- 0x1c9e
		"01011010",	-- 0x1c9f
		"00010100",	-- 0x1ca0
		"00110101",	-- 0x1ca1
		"00011111",	-- 0x1ca2
		"00010001",	-- 0x1ca3
		"00110111",	-- 0x1ca4
		"01010110",	-- 0x1ca5
		"00001110",	-- 0x1ca6
		"00110111",	-- 0x1ca7
		"10011001",	-- 0x1ca8
		"00001011",	-- 0x1ca9
		"01111001",	-- 0x1caa
		"00001010",	-- 0x1cab
		"01011101",	-- 0x1cac
		"01000101",	-- 0x1cad
		"00000110",	-- 0x1cae
		"11001100",	-- 0x1caf
		"00011000",	-- 0x1cb0
		"01000100",	-- 0x1cb1
		"00000010",	-- 0x1cb2
		"01110010",	-- 0x1cb3
		"10110110",	-- 0x1cb4
		"11011010",	-- 0x1cb5
		"01001111",	-- 0x1cb6
		"10110010",	-- 0x1cb7
		"00000001",	-- 0x1cb8
		"11011010",	-- 0x1cb9
		"11111010",	-- 0x1cba
		"00000001",	-- 0x1cbb
		"11011011",	-- 0x1cbc
		"10010010",	-- 0x1cbd
		"01001111",	-- 0x1cbe
		"01111001",	-- 0x1cbf
		"00110100",	-- 0x1cc0
		"01011001",	-- 0x1cc1
		"01000100",	-- 0x1cc2
		"00000010",	-- 0x1cc3
		"01110101",	-- 0x1cc4
		"00011111",	-- 0x1cc5
		"01111001",	-- 0x1cc6
		"00111100",	-- 0x1cc7
		"01011001",	-- 0x1cc8
		"01000101",	-- 0x1cc9
		"00000010",	-- 0x1cca
		"01110111",	-- 0x1ccb
		"00011111",	-- 0x1ccc
		"11011010",	-- 0x1ccd
		"11001010",	-- 0x1cce
		"00110111",	-- 0x1ccf
		"10011010",	-- 0x1cd0
		"00000110",	-- 0x1cd1
		"00110111",	-- 0x1cd2
		"10111010",	-- 0x1cd3
		"00001010",	-- 0x1cd4
		"00110111",	-- 0x1cd5
		"00111001",	-- 0x1cd6
		"00000111",	-- 0x1cd7
		"11001100",	-- 0x1cd8
		"00011000",	-- 0x1cd9
		"01000100",	-- 0x1cda
		"00000011",	-- 0x1cdb
		"01010010",	-- 0x1cdc
		"10010010",	-- 0x1cdd
		"11001010",	-- 0x1cde
		"11111011",	-- 0x1cdf
		"00000001",	-- 0x1ce0
		"11011100",	-- 0x1ce1
		"11001111",	-- 0x1ce2
		"00000100",	-- 0x1ce3
		"01000110",	-- 0x1ce4
		"00011100",	-- 0x1ce5
		"11011010",	-- 0x1ce6
		"11001010",	-- 0x1ce7
		"11001100",	-- 0x1ce8
		"00011000",	-- 0x1ce9
		"01000100",	-- 0x1cea
		"00010110",	-- 0x1ceb
		"00110111",	-- 0x1cec
		"00111001",	-- 0x1ced
		"00010011",	-- 0x1cee
		"00110111",	-- 0x1cef
		"10011010",	-- 0x1cf0
		"00010000",	-- 0x1cf1
		"00110111",	-- 0x1cf2
		"10111010",	-- 0x1cf3
		"00001101",	-- 0x1cf4
		"00110101",	-- 0x1cf5
		"10011001",	-- 0x1cf6
		"00001010",	-- 0x1cf7
		"01111001",	-- 0x1cf8
		"00011001",	-- 0x1cf9
		"01011101",	-- 0x1cfa
		"01000101",	-- 0x1cfb
		"00000101",	-- 0x1cfc
		"00110101",	-- 0x1cfd
		"00011111",	-- 0x1cfe
		"00000010",	-- 0x1cff
		"01110010",	-- 0x1d00
		"10110111",	-- 0x1d01
		"11011010",	-- 0x1d02
		"01001111",	-- 0x1d03
		"10110010",	-- 0x1d04
		"00000001",	-- 0x1d05
		"11011011",	-- 0x1d06
		"01010010",	-- 0x1d07
		"10110010",	-- 0x1d08
		"00000001",	-- 0x1d09
		"01101000",	-- 0x1d0a
		"11111010",	-- 0x1d0b
		"00000001",	-- 0x1d0c
		"11001111",	-- 0x1d0d
		"10010010",	-- 0x1d0e
		"01001110",	-- 0x1d0f
		"01111001",	-- 0x1d10
		"10001101",	-- 0x1d11
		"01010110",	-- 0x1d12
		"01000010",	-- 0x1d13
		"00000010",	-- 0x1d14
		"01110111",	-- 0x1d15
		"00011110",	-- 0x1d16
		"00110101",	-- 0x1d17
		"00011001",	-- 0x1d18
		"00000100",	-- 0x1d19
		"01110101",	-- 0x1d1a
		"00011110",	-- 0x1d1b
		"01110010",	-- 0x1d1c
		"11100101",	-- 0x1d1d
		"01111001",	-- 0x1d1e
		"00011111",	-- 0x1d1f
		"11100101",	-- 0x1d20
		"01000101",	-- 0x1d21
		"00000101",	-- 0x1d22
		"00110111",	-- 0x1d23
		"00011110",	-- 0x1d24
		"00000010",	-- 0x1d25
		"01110111",	-- 0x1d26
		"00011011",	-- 0x1d27
		"01000000",	-- 0x1d28
		"00001110",	-- 0x1d29
		"00110101",	-- 0x1d2a
		"01010000",	-- 0x1d2b
		"00000010",	-- 0x1d2c
		"01110101",	-- 0x1d2d
		"00111011",	-- 0x1d2e
		"11011011",	-- 0x1d2f
		"10100010",	-- 0x1d30
		"01001011",	-- 0x1d31
		"00000100",	-- 0x1d32
		"01110010",	-- 0x1d33
		"11100101",	-- 0x1d34
		"01110101",	-- 0x1d35
		"00011011",	-- 0x1d36
		"01100011",	-- 0x1d37
		"11011010",	-- 0x1d38
		"01001110",	-- 0x1d39
		"10110010",	-- 0x1d3a
		"00000001",	-- 0x1d3b
		"11001111",	-- 0x1d3c
		"00110111",	-- 0x1d3d
		"00011001",	-- 0x1d3e
		"00000010",	-- 0x1d3f
		"01110101",	-- 0x1d40
		"11111101",	-- 0x1d41
		"01111001",	-- 0x1d42
		"00010100",	-- 0x1d43
		"01011001",	-- 0x1d44
		"01000101",	-- 0x1d45
		"00001010",	-- 0x1d46
		"01111001",	-- 0x1d47
		"00000111",	-- 0x1d48
		"11000111",	-- 0x1d49
		"01000101",	-- 0x1d4a
		"00000101",	-- 0x1d4b
		"00110111",	-- 0x1d4c
		"11111101",	-- 0x1d4d
		"00000010",	-- 0x1d4e
		"01110111",	-- 0x1d4f
		"00111011",	-- 0x1d50
		"01000000",	-- 0x1d51
		"00000110",	-- 0x1d52
		"00110101",	-- 0x1d53
		"00011001",	-- 0x1d54
		"00000010",	-- 0x1d55
		"01110111",	-- 0x1d56
		"11111101",	-- 0x1d57
		"01100011",	-- 0x1d58
		"00110111",	-- 0x1d59
		"00100000",	-- 0x1d5a
		"00001000",	-- 0x1d5b
		"00110101",	-- 0x1d5c
		"11011101",	-- 0x1d5d
		"00000111",	-- 0x1d5e
		"01110111",	-- 0x1d5f
		"11011101",	-- 0x1d60
		"01110010",	-- 0x1d61
		"11000010",	-- 0x1d62
		"10001100",	-- 0x1d63
		"01110101",	-- 0x1d64
		"11011101",	-- 0x1d65
		"00000011",	-- 0x1d66
		"11100001",	-- 0x1d67
		"00010010",	-- 0x1d68
		"11111010",	-- 0x1d69
		"00000010",	-- 0x1d6a
		"01000010",	-- 0x1d6b
		"11001110",	-- 0x1d6c
		"00001000",	-- 0x1d6d
		"01000111",	-- 0x1d6e
		"00000011",	-- 0x1d6f
		"01110111",	-- 0x1d70
		"11111100",	-- 0x1d71
		"10001100",	-- 0x1d72
		"01110101",	-- 0x1d73
		"11111100",	-- 0x1d74
		"11001110",	-- 0x1d75
		"00010000",	-- 0x1d76
		"01000111",	-- 0x1d77
		"00000011",	-- 0x1d78
		"01110111",	-- 0x1d79
		"01011100",	-- 0x1d7a
		"10001100",	-- 0x1d7b
		"01110101",	-- 0x1d7c
		"01011100",	-- 0x1d7d
		"00110101",	-- 0x1d7e
		"11011001",	-- 0x1d7f
		"00011111",	-- 0x1d80
		"00110111",	-- 0x1d81
		"01010000",	-- 0x1d82
		"00010010",	-- 0x1d83
		"01110101",	-- 0x1d84
		"01010000",	-- 0x1d85
		"00110101",	-- 0x1d86
		"01111000",	-- 0x1d87
		"00000011",	-- 0x1d88
		"00110111",	-- 0x1d89
		"00111101",	-- 0x1d8a
		"00001010",	-- 0x1d8b
		"01110101",	-- 0x1d8c
		"00111101",	-- 0x1d8d
		"10010110",	-- 0x1d8e
		"01001011",	-- 0x1d8f
		"11000010",	-- 0x1d90
		"11000101",	-- 0x1d91
		"11000011",	-- 0x1d92
		"00000101",	-- 0x1d93
		"10011010",	-- 0x1d94
		"01001011",	-- 0x1d95
		"01110101",	-- 0x1d96
		"01111000",	-- 0x1d97
		"11011010",	-- 0x1d98
		"10100000",	-- 0x1d99
		"11000010",	-- 0x1d9a
		"01110000",	-- 0x1d9b
		"10010010",	-- 0x1d9c
		"10100000",	-- 0x1d9d
		"01110101",	-- 0x1d9e
		"10111000",	-- 0x1d9f
		"00110111",	-- 0x1da0
		"11011001",	-- 0x1da1
		"00010101",	-- 0x1da2
		"10110110",	-- 0x1da3
		"00000001",	-- 0x1da4
		"00001010",	-- 0x1da5
		"10110111",	-- 0x1da6
		"00000001",	-- 0x1da7
		"00011010",	-- 0x1da8
		"00000001",	-- 0x1da9
		"11000100",	-- 0x1daa
		"11011100",	-- 0x1dab
		"10110011",	-- 0x1dac
		"00000010",	-- 0x1dad
		"00010111",	-- 0x1dae
		"10110110",	-- 0x1daf
		"00000001",	-- 0x1db0
		"10011000",	-- 0x1db1
		"00000001",	-- 0x1db2
		"11000100",	-- 0x1db3
		"11011111",	-- 0x1db4
		"10110011",	-- 0x1db5
		"00000010",	-- 0x1db6
		"00011001",	-- 0x1db7
		"11111010",	-- 0x1db8
		"00000001",	-- 0x1db9
		"11001111",	-- 0x1dba
		"10010010",	-- 0x1dbb
		"01001110",	-- 0x1dbc
		"11111010",	-- 0x1dbd
		"00000001",	-- 0x1dbe
		"11011001",	-- 0x1dbf
		"10010010",	-- 0x1dc0
		"01001111",	-- 0x1dc1
		"00110111",	-- 0x1dc2
		"01011111",	-- 0x1dc3
		"01000011",	-- 0x1dc4
		"01111001",	-- 0x1dc5
		"00011110",	-- 0x1dc6
		"01011001",	-- 0x1dc7
		"01000101",	-- 0x1dc8
		"00111110",	-- 0x1dc9
		"01111001",	-- 0x1dca
		"01100100",	-- 0x1dcb
		"01011101",	-- 0x1dcc
		"01000100",	-- 0x1dcd
		"00111001",	-- 0x1dce
		"01111001",	-- 0x1dcf
		"00101101",	-- 0x1dd0
		"01010000",	-- 0x1dd1
		"01000101",	-- 0x1dd2
		"00110100",	-- 0x1dd3
		"11011011",	-- 0x1dd4
		"10000100",	-- 0x1dd5
		"11001111",	-- 0x1dd6
		"01000000",	-- 0x1dd7
		"01000110",	-- 0x1dd8
		"00101110",	-- 0x1dd9
		"11011011",	-- 0x1dda
		"10000000",	-- 0x1ddb
		"11001111",	-- 0x1ddc
		"00001000",	-- 0x1ddd
		"01000110",	-- 0x1dde
		"00101000",	-- 0x1ddf
		"11011011",	-- 0x1de0
		"10000000",	-- 0x1de1
		"11001111",	-- 0x1de2
		"01000000",	-- 0x1de3
		"01000110",	-- 0x1de4
		"00100010",	-- 0x1de5
		"11011011",	-- 0x1de6
		"10000000",	-- 0x1de7
		"11001111",	-- 0x1de8
		"00100000",	-- 0x1de9
		"01000110",	-- 0x1dea
		"00011100",	-- 0x1deb
		"11011011",	-- 0x1dec
		"10000010",	-- 0x1ded
		"11001111",	-- 0x1dee
		"01000000",	-- 0x1def
		"01000110",	-- 0x1df0
		"00010110",	-- 0x1df1
		"00110111",	-- 0x1df2
		"11111111",	-- 0x1df3
		"00010011",	-- 0x1df4
		"10111110",	-- 0x1df5
		"00000001",	-- 0x1df6
		"10000111",	-- 0x1df7
		"10001100",	-- 0x1df8
		"00000001",	-- 0x1df9
		"00110001",	-- 0x1dfa
		"01000100",	-- 0x1dfb
		"00001011",	-- 0x1dfc
		"11111010",	-- 0x1dfd
		"00000001",	-- 0x1dfe
		"10000110",	-- 0x1dff
		"11001100",	-- 0x1e00
		"01001000",	-- 0x1e01
		"01000101",	-- 0x1e02
		"00000100",	-- 0x1e03
		"11001100",	-- 0x1e04
		"10001111",	-- 0x1e05
		"01000101",	-- 0x1e06
		"00000010",	-- 0x1e07
		"01110010",	-- 0x1e08
		"11101100",	-- 0x1e09
		"01111001",	-- 0x1e0a
		"00111100",	-- 0x1e0b
		"11101100",	-- 0x1e0c
		"01000101",	-- 0x1e0d
		"00001101",	-- 0x1e0e
		"01110111",	-- 0x1e0f
		"10111100",	-- 0x1e10
		"00110111",	-- 0x1e11
		"01010000",	-- 0x1e12
		"00001000",	-- 0x1e13
		"11011011",	-- 0x1e14
		"10100000",	-- 0x1e15
		"11000111",	-- 0x1e16
		"00100000",	-- 0x1e17
		"10010011",	-- 0x1e18
		"10100000",	-- 0x1e19
		"01110111",	-- 0x1e1a
		"01111000",	-- 0x1e1b
		"00110111",	-- 0x1e1c
		"00110110",	-- 0x1e1d
		"00110001",	-- 0x1e1e
		"11111011",	-- 0x1e1f
		"00000001",	-- 0x1e20
		"10000101",	-- 0x1e21
		"01111001",	-- 0x1e22
		"00001010",	-- 0x1e23
		"11101101",	-- 0x1e24
		"01000100",	-- 0x1e25
		"00011011",	-- 0x1e26
		"11111010",	-- 0x1e27
		"00000001",	-- 0x1e28
		"10000110",	-- 0x1e29
		"11001100",	-- 0x1e2a
		"01001000",	-- 0x1e2b
		"01000100",	-- 0x1e2c
		"00000010",	-- 0x1e2d
		"01110111",	-- 0x1e2e
		"00111110",	-- 0x1e2f
		"11001100",	-- 0x1e30
		"10001111",	-- 0x1e31
		"01000101",	-- 0x1e32
		"00100100",	-- 0x1e33
		"00110111",	-- 0x1e34
		"00111110",	-- 0x1e35
		"00100001",	-- 0x1e36
		"01010111",	-- 0x1e37
		"01000110",	-- 0x1e38
		"00000001",	-- 0x1e39
		"01010001",	-- 0x1e3a
		"10110011",	-- 0x1e3b
		"00000001",	-- 0x1e3c
		"10000101",	-- 0x1e3d
		"01110101",	-- 0x1e3e
		"00111110",	-- 0x1e3f
		"01000000",	-- 0x1e40
		"00010110",	-- 0x1e41
		"11001101",	-- 0x1e42
		"00000100",	-- 0x1e43
		"01000101",	-- 0x1e44
		"00001010",	-- 0x1e45
		"00110101",	-- 0x1e46
		"01010000",	-- 0x1e47
		"00000111",	-- 0x1e48
		"11001010",	-- 0x1e49
		"11011111",	-- 0x1e4a
		"00000001",	-- 0x1e4b
		"11011111",	-- 0x1e4c
		"10101010",	-- 0x1e4d
		"01110101",	-- 0x1e4e
		"10111100",	-- 0x1e4f
		"01010011",	-- 0x1e50
		"10110011",	-- 0x1e51
		"00000001",	-- 0x1e52
		"10000101",	-- 0x1e53
		"01110101",	-- 0x1e54
		"00111110",	-- 0x1e55
		"01110010",	-- 0x1e56
		"11101101",	-- 0x1e57
		"01000000",	-- 0x1e58
		"00100001",	-- 0x1e59
		"01110101",	-- 0x1e5a
		"11111111",	-- 0x1e5b
		"10111110",	-- 0x1e5c
		"00000001",	-- 0x1e5d
		"10000111",	-- 0x1e5e
		"10001100",	-- 0x1e5f
		"00000000",	-- 0x1e60
		"00000011",	-- 0x1e61
		"01000101",	-- 0x1e62
		"00000111",	-- 0x1e63
		"10001100",	-- 0x1e64
		"00000001",	-- 0x1e65
		"00110001",	-- 0x1e66
		"01000100",	-- 0x1e67
		"00000010",	-- 0x1e68
		"01110111",	-- 0x1e69
		"11111111",	-- 0x1e6a
		"01010010",	-- 0x1e6b
		"01010011",	-- 0x1e6c
		"10111010",	-- 0x1e6d
		"00000001",	-- 0x1e6e
		"10000111",	-- 0x1e6f
		"01100011",	-- 0x1e70
		"10111110",	-- 0x1e71
		"00000001",	-- 0x1e72
		"10000111",	-- 0x1e73
		"00011100",	-- 0x1e74
		"01000111",	-- 0x1e75
		"00000011",	-- 0x1e76
		"00001010",	-- 0x1e77
		"00000001",	-- 0x1e78
		"10000111",	-- 0x1e79
		"01100011",	-- 0x1e7a
		"11011010",	-- 0x1e7b
		"01001110",	-- 0x1e7c
		"10110010",	-- 0x1e7d
		"00000001",	-- 0x1e7e
		"11001111",	-- 0x1e7f
		"00110101",	-- 0x1e80
		"11010000",	-- 0x1e81
		"00111110",	-- 0x1e82
		"11011010",	-- 0x1e83
		"01011101",	-- 0x1e84
		"01000110",	-- 0x1e85
		"00100100",	-- 0x1e86
		"01111001",	-- 0x1e87
		"00101000",	-- 0x1e88
		"01011001",	-- 0x1e89
		"01000101",	-- 0x1e8a
		"00100001",	-- 0x1e8b
		"01111001",	-- 0x1e8c
		"01100100",	-- 0x1e8d
		"01011001",	-- 0x1e8e
		"01000100",	-- 0x1e8f
		"00011100",	-- 0x1e90
		"01111001",	-- 0x1e91
		"00110011",	-- 0x1e92
		"01010000",	-- 0x1e93
		"01000101",	-- 0x1e94
		"00010111",	-- 0x1e95
		"01111001",	-- 0x1e96
		"11100100",	-- 0x1e97
		"01010111",	-- 0x1e98
		"01000011",	-- 0x1e99
		"00010010",	-- 0x1e9a
		"00110101",	-- 0x1e9b
		"11010011",	-- 0x1e9c
		"00001111",	-- 0x1e9d
		"11011010",	-- 0x1e9e
		"10000000",	-- 0x1e9f
		"11001110",	-- 0x1ea0
		"00001000",	-- 0x1ea1
		"01000110",	-- 0x1ea2
		"00001001",	-- 0x1ea3
		"11011010",	-- 0x1ea4
		"10000000",	-- 0x1ea5
		"11001110",	-- 0x1ea6
		"00100000",	-- 0x1ea7
		"01000111",	-- 0x1ea8
		"00000101",	-- 0x1ea9
		"10001100",	-- 0x1eaa
		"01110101",	-- 0x1eab
		"11011011",	-- 0x1eac
		"01110010",	-- 0x1ead
		"11100110",	-- 0x1eae
		"01111001",	-- 0x1eaf
		"01111010",	-- 0x1eb0
		"11100110",	-- 0x1eb1
		"01000101",	-- 0x1eb2
		"00000010",	-- 0x1eb3
		"01110111",	-- 0x1eb4
		"11011011",	-- 0x1eb5
		"01111001",	-- 0x1eb6
		"00000101",	-- 0x1eb7
		"01011101",	-- 0x1eb8
		"01000101",	-- 0x1eb9
		"00000110",	-- 0x1eba
		"11011010",	-- 0x1ebb
		"10100000",	-- 0x1ebc
		"11000010",	-- 0x1ebd
		"11111011",	-- 0x1ebe
		"10010010",	-- 0x1ebf
		"10100000",	-- 0x1ec0
		"00110111",	-- 0x1ec1
		"10111111",	-- 0x1ec2
		"00011111",	-- 0x1ec3
		"01111001",	-- 0x1ec4
		"00011110",	-- 0x1ec5
		"01011001",	-- 0x1ec6
		"01000101",	-- 0x1ec7
		"00011010",	-- 0x1ec8
		"01111001",	-- 0x1ec9
		"01100100",	-- 0x1eca
		"01011101",	-- 0x1ecb
		"01000100",	-- 0x1ecc
		"00010101",	-- 0x1ecd
		"01111001",	-- 0x1ece
		"11011100",	-- 0x1ecf
		"01010111",	-- 0x1ed0
		"01000101",	-- 0x1ed1
		"00010000",	-- 0x1ed2
		"11011010",	-- 0x1ed3
		"10000000",	-- 0x1ed4
		"11001110",	-- 0x1ed5
		"01000000",	-- 0x1ed6
		"01000110",	-- 0x1ed7
		"00001010",	-- 0x1ed8
		"11011010",	-- 0x1ed9
		"10000000",	-- 0x1eda
		"11001110",	-- 0x1edb
		"00001000",	-- 0x1edc
		"01000110",	-- 0x1edd
		"00000100",	-- 0x1ede
		"11011010",	-- 0x1edf
		"01011111",	-- 0x1ee0
		"01001010",	-- 0x1ee1
		"00000010",	-- 0x1ee2
		"01110010",	-- 0x1ee3
		"11101110",	-- 0x1ee4
		"01111001",	-- 0x1ee5
		"01011010",	-- 0x1ee6
		"11101110",	-- 0x1ee7
		"01000101",	-- 0x1ee8
		"00001101",	-- 0x1ee9
		"01110111",	-- 0x1eea
		"11011100",	-- 0x1eeb
		"00110111",	-- 0x1eec
		"01010000",	-- 0x1eed
		"00001000",	-- 0x1eee
		"11011010",	-- 0x1eef
		"10100000",	-- 0x1ef0
		"11000110",	-- 0x1ef1
		"01000000",	-- 0x1ef2
		"10010010",	-- 0x1ef3
		"10100000",	-- 0x1ef4
		"01110111",	-- 0x1ef5
		"01111000",	-- 0x1ef6
		"11011010",	-- 0x1ef7
		"01011111",	-- 0x1ef8
		"01001010",	-- 0x1ef9
		"00001010",	-- 0x1efa
		"00110101",	-- 0x1efb
		"01010000",	-- 0x1efc
		"00000111",	-- 0x1efd
		"01110101",	-- 0x1efe
		"11011100",	-- 0x1eff
		"11001010",	-- 0x1f00
		"10111111",	-- 0x1f01
		"00000001",	-- 0x1f02
		"11011111",	-- 0x1f03
		"10101010",	-- 0x1f04
		"00110111",	-- 0x1f05
		"01010000",	-- 0x1f06
		"00010111",	-- 0x1f07
		"00110111",	-- 0x1f08
		"10111001",	-- 0x1f09
		"00010100",	-- 0x1f0a
		"00110101",	-- 0x1f0b
		"00011001",	-- 0x1f0c
		"00010001",	-- 0x1f0d
		"01111001",	-- 0x1f0e
		"01011100",	-- 0x1f0f
		"11010000",	-- 0x1f10
		"01000101",	-- 0x1f11
		"00000011",	-- 0x1f12
		"00110111",	-- 0x1f13
		"00111001",	-- 0x1f14
		"00000110",	-- 0x1f15
		"00110101",	-- 0x1f16
		"01111001",	-- 0x1f17
		"00000011",	-- 0x1f18
		"00110101",	-- 0x1f19
		"11010010",	-- 0x1f1a
		"00000011",	-- 0x1f1b
		"01110111",	-- 0x1f1c
		"10111000",	-- 0x1f1d
		"10001100",	-- 0x1f1e
		"01110101",	-- 0x1f1f
		"10111000",	-- 0x1f20
		"00110111",	-- 0x1f21
		"00011001",	-- 0x1f22
		"00000110",	-- 0x1f23
		"11011010",	-- 0x1f24
		"10100000",	-- 0x1f25
		"11000010",	-- 0x1f26
		"11110111",	-- 0x1f27
		"10010010",	-- 0x1f28
		"10100000",	-- 0x1f29
		"11111010",	-- 0x1f2a
		"00000001",	-- 0x1f2b
		"11010101",	-- 0x1f2c
		"10010010",	-- 0x1f2d
		"01001110",	-- 0x1f2e
		"00000101",	-- 0x1f2f
		"10010110",	-- 0x1f30
		"01001011",	-- 0x1f31
		"00110111",	-- 0x1f32
		"10101010",	-- 0x1f33
		"00000101",	-- 0x1f34
		"01111001",	-- 0x1f35
		"01111010",	-- 0x1f36
		"10111111",	-- 0x1f37
		"01000010",	-- 0x1f38
		"00000101",	-- 0x1f39
		"01110101",	-- 0x1f3a
		"10011101",	-- 0x1f3b
		"01010010",	-- 0x1f3c
		"01000000",	-- 0x1f3d
		"00100001",	-- 0x1f3e
		"00110101",	-- 0x1f3f
		"10101101",	-- 0x1f40
		"00010000",	-- 0x1f41
		"00110101",	-- 0x1f42
		"10101001",	-- 0x1f43
		"00001101",	-- 0x1f44
		"01111001",	-- 0x1f45
		"01111010",	-- 0x1f46
		"10111110",	-- 0x1f47
		"01000011",	-- 0x1f48
		"00001000",	-- 0x1f49
		"00110101",	-- 0x1f4a
		"00011001",	-- 0x1f4b
		"00000101",	-- 0x1f4c
		"01111001",	-- 0x1f4d
		"01111010",	-- 0x1f4e
		"11000000",	-- 0x1f4f
		"01000010",	-- 0x1f50
		"00010100",	-- 0x1f51
		"11000010",	-- 0x1f52
		"10000101",	-- 0x1f53
		"01110101",	-- 0x1f54
		"11111110",	-- 0x1f55
		"01110101",	-- 0x1f56
		"10011000",	-- 0x1f57
		"01101100",	-- 0x1f58
		"11011010",	-- 0x1f59
		"01101101",	-- 0x1f5a
		"11000010",	-- 0x1f5b
		"11111110",	-- 0x1f5c
		"10010010",	-- 0x1f5d
		"01101101",	-- 0x1f5e
		"01111100",	-- 0x1f5f
		"11000011",	-- 0x1f60
		"00000001",	-- 0x1f61
		"10011010",	-- 0x1f62
		"01001011",	-- 0x1f63
		"01110101",	-- 0x1f64
		"01111000",	-- 0x1f65
		"10011010",	-- 0x1f66
		"01111000",	-- 0x1f67
		"00110111",	-- 0x1f68
		"01111000",	-- 0x1f69
		"00000010",	-- 0x1f6a
		"01110111",	-- 0x1f6b
		"00111101",	-- 0x1f6c
		"00000111",	-- 0x1f6d
		"00000001",	-- 0x1f6e
		"11110111",	-- 0x1f6f
		"01100001",	-- 0x1f70
		"01101100",	-- 0x1f71
		"01011010",	-- 0x1f72
		"11000011",	-- 0x1f73
		"00011111",	-- 0x1f74
		"10001110",	-- 0x1f75
		"00000000",	-- 0x1f76
		"10000010",	-- 0x1f77
		"11100111",	-- 0x1f78
		"00000000",	-- 0x1f79
		"11010010",	-- 0x1f7a
		"10100000",	-- 0x1f7b
		"11000010",	-- 0x1f7c
		"01100000",	-- 0x1f7d
		"10010010",	-- 0x1f7e
		"01111010",	-- 0x1f7f
		"11010111",	-- 0x1f80
		"01111010",	-- 0x1f81
		"00000001",	-- 0x1f82
		"11010001",	-- 0x1f83
		"10011000",	-- 0x1f84
		"01111101",	-- 0x1f85
		"11000011",	-- 0x1f86
		"11111111",	-- 0x1f87
		"10001110",	-- 0x1f88
		"00000000",	-- 0x1f89
		"10000000",	-- 0x1f8a
		"11100111",	-- 0x1f8b
		"00000000",	-- 0x1f8c
		"00000001",	-- 0x1f8d
		"11010001",	-- 0x1f8e
		"10011000",	-- 0x1f8f
		"11011011",	-- 0x1f90
		"01111001",	-- 0x1f91
		"11000011",	-- 0x1f92
		"01100000",	-- 0x1f93
		"11010111",	-- 0x1f94
		"10000100",	-- 0x1f95
		"00110111",	-- 0x1f96
		"11111110",	-- 0x1f97
		"00000010",	-- 0x1f98
		"11000111",	-- 0x1f99
		"00000001",	-- 0x1f9a
		"10001110",	-- 0x1f9b
		"00000000",	-- 0x1f9c
		"10000100",	-- 0x1f9d
		"00000001",	-- 0x1f9e
		"11010001",	-- 0x1f9f
		"10011000",	-- 0x1fa0
		"01000000",	-- 0x1fa1
		"00010101",	-- 0x1fa2
		"11011010",	-- 0x1fa3
		"10000100",	-- 0x1fa4
		"11000010",	-- 0x1fa5
		"01100000",	-- 0x1fa6
		"10010010",	-- 0x1fa7
		"10100000",	-- 0x1fa8
		"01100011",	-- 0x1fa9
		"01011011",	-- 0x1faa
		"11010010",	-- 0x1fab
		"10100000",	-- 0x1fac
		"10010010",	-- 0x1fad
		"10100000",	-- 0x1fae
		"10001110",	-- 0x1faf
		"00000000",	-- 0x1fb0
		"10000100",	-- 0x1fb1
		"11100011",	-- 0x1fb2
		"00000000",	-- 0x1fb3
		"00000001",	-- 0x1fb4
		"11010001",	-- 0x1fb5
		"10011000",	-- 0x1fb6
		"01100011",	-- 0x1fb7
		"11011010",	-- 0x1fb8
		"01001110",	-- 0x1fb9
		"10110010",	-- 0x1fba
		"00000001",	-- 0x1fbb
		"11010101",	-- 0x1fbc
		"01010010",	-- 0x1fbd
		"00000001",	-- 0x1fbe
		"11100000",	-- 0x1fbf
		"10100101",	-- 0x1fc0
		"01000111",	-- 0x1fc1
		"00000011",	-- 0x1fc2
		"01110111",	-- 0x1fc3
		"10010110",	-- 0x1fc4
		"10001100",	-- 0x1fc5
		"01110101",	-- 0x1fc6
		"10010110",	-- 0x1fc7
		"00110101",	-- 0x1fc8
		"10101010",	-- 0x1fc9
		"00000011",	-- 0x1fca
		"00000011",	-- 0x1fcb
		"11100000",	-- 0x1fcc
		"10001101",	-- 0x1fcd
		"00110101",	-- 0x1fce
		"10111001",	-- 0x1fcf
		"00000011",	-- 0x1fd0
		"00110111",	-- 0x1fd1
		"00011101",	-- 0x1fd2
		"01101010",	-- 0x1fd3
		"11011010",	-- 0x1fd4
		"10101001",	-- 0x1fd5
		"01010110",	-- 0x1fd6
		"01000111",	-- 0x1fd7
		"00100110",	-- 0x1fd8
		"11111011",	-- 0x1fd9
		"00000001",	-- 0x1fda
		"10000011",	-- 0x1fdb
		"01010111",	-- 0x1fdc
		"01000110",	-- 0x1fdd
		"00101110",	-- 0x1fde
		"11011010",	-- 0x1fdf
		"10101000",	-- 0x1fe0
		"01000111",	-- 0x1fe1
		"00011100",	-- 0x1fe2
		"01010000",	-- 0x1fe3
		"01000111",	-- 0x1fe4
		"00001100",	-- 0x1fe5
		"11001011",	-- 0x1fe6
		"01111000",	-- 0x1fe7
		"11001110",	-- 0x1fe8
		"00001111",	-- 0x1fe9
		"01000110",	-- 0x1fea
		"01001110",	-- 0x1feb
		"10000001",	-- 0x1fec
		"00010000",	-- 0x1fed
		"11001011",	-- 0x1fee
		"01101001",	-- 0x1fef
		"01000000",	-- 0x1ff0
		"01001000",	-- 0x1ff1
		"10010010",	-- 0x1ff2
		"10101000",	-- 0x1ff3
		"11011010",	-- 0x1ff4
		"10101001",	-- 0x1ff5
		"00000001",	-- 0x1ff6
		"11100000",	-- 0x1ff7
		"10100101",	-- 0x1ff8
		"01000111",	-- 0x1ff9
		"00001101",	-- 0x1ffa
		"11001011",	-- 0x1ffb
		"01011010",	-- 0x1ffc
		"01000000",	-- 0x1ffd
		"00101101",	-- 0x1ffe
		"00000001",	-- 0x1fff
		"11100000",	-- 0x2000
		"10100101",	-- 0x2001
		"01000110",	-- 0x2002
		"00000100",	-- 0x2003
		"11001011",	-- 0x2004
		"01111100",	-- 0x2005
		"01000000",	-- 0x2006
		"00100010",	-- 0x2007
		"01010010",	-- 0x2008
		"11001011",	-- 0x2009
		"00111011",	-- 0x200a
		"01000000",	-- 0x200b
		"00011111",	-- 0x200c
		"01001001",	-- 0x200d
		"00000011",	-- 0x200e
		"00000011",	-- 0x200f
		"11100000",	-- 0x2010
		"10011001",	-- 0x2011
		"11011010",	-- 0x2012
		"10101000",	-- 0x2013
		"01000110",	-- 0x2014
		"00100010",	-- 0x2015
		"10110010",	-- 0x2016
		"00000001",	-- 0x2017
		"10000011",	-- 0x2018
		"00110111",	-- 0x2019
		"10111001",	-- 0x201a
		"00100010",	-- 0x201b
		"01110111",	-- 0x201c
		"00011101",	-- 0x201d
		"11011010",	-- 0x201e
		"10101001",	-- 0x201f
		"01001011",	-- 0x2020
		"00000110",	-- 0x2021
		"01000110",	-- 0x2022
		"00001100",	-- 0x2023
		"01100001",	-- 0x2024
		"01111111",	-- 0x2025
		"01000110",	-- 0x2026
		"00001000",	-- 0x2027
		"11001011",	-- 0x2028
		"11111100",	-- 0x2029
		"11001010",	-- 0x202a
		"10000000",	-- 0x202b
		"10010010",	-- 0x202c
		"10101001",	-- 0x202d
		"01000000",	-- 0x202e
		"01101001",	-- 0x202f
		"10010010",	-- 0x2030
		"10101001",	-- 0x2031
		"10001111",	-- 0x2032
		"11100000",	-- 0x2033
		"11001100",	-- 0x2034
		"00001101",	-- 0x2035
		"11101010",	-- 0x2036
		"10000010",	-- 0x2037
		"11001011",	-- 0x2038
		"11111000",	-- 0x2039
		"10010010",	-- 0x203a
		"10101000",	-- 0x203b
		"01000000",	-- 0x203c
		"01011011",	-- 0x203d
		"00110111",	-- 0x203e
		"01010000",	-- 0x203f
		"00011110",	-- 0x2040
		"00110111",	-- 0x2041
		"00010110",	-- 0x2042
		"00011011",	-- 0x2043
		"11111011",	-- 0x2044
		"00000001",	-- 0x2045
		"10000011",	-- 0x2046
		"11001101",	-- 0x2047
		"01111110",	-- 0x2048
		"01000100",	-- 0x2049
		"00000010",	-- 0x204a
		"11001011",	-- 0x204b
		"01111111",	-- 0x204c
		"11001101",	-- 0x204d
		"11111110",	-- 0x204e
		"01001100",	-- 0x204f
		"00000010",	-- 0x2050
		"11001011",	-- 0x2051
		"11111111",	-- 0x2052
		"01010111",	-- 0x2053
		"01000111",	-- 0x2054
		"00000101",	-- 0x2055
		"01001000",	-- 0x2056
		"00000101",	-- 0x2057
		"11001011",	-- 0x2058
		"11111110",	-- 0x2059
		"10001100",	-- 0x205a
		"11001011",	-- 0x205b
		"01111110",	-- 0x205c
		"01000000",	-- 0x205d
		"00110011",	-- 0x205e
		"00110111",	-- 0x205f
		"01010000",	-- 0x2060
		"00000101",	-- 0x2061
		"11001011",	-- 0x2062
		"11111110",	-- 0x2063
		"00110101",	-- 0x2064
		"00111101",	-- 0x2065
		"00101011",	-- 0x2066
		"11001011",	-- 0x2067
		"10110100",	-- 0x2068
		"11011010",	-- 0x2069
		"01111000",	-- 0x206a
		"11000010",	-- 0x206b
		"11101111",	-- 0x206c
		"01000110",	-- 0x206d
		"00100011",	-- 0x206e
		"11011010",	-- 0x206f
		"01111001",	-- 0x2070
		"11000010",	-- 0x2071
		"00000001",	-- 0x2072
		"01000110",	-- 0x2073
		"00011101",	-- 0x2074
		"11111010",	-- 0x2075
		"00000001",	-- 0x2076
		"11010101",	-- 0x2077
		"11001110",	-- 0x2078
		"10000000",	-- 0x2079
		"01000110",	-- 0x207a
		"00010110",	-- 0x207b
		"11011010",	-- 0x207c
		"01101101",	-- 0x207d
		"11001110",	-- 0x207e
		"00000001",	-- 0x207f
		"01000110",	-- 0x2080
		"00010000",	-- 0x2081
		"00110101",	-- 0x2082
		"10011000",	-- 0x2083
		"00001101",	-- 0x2084
		"11111011",	-- 0x2085
		"00000001",	-- 0x2086
		"10000011",	-- 0x2087
		"01010111",	-- 0x2088
		"01001010",	-- 0x2089
		"00000010",	-- 0x208a
		"01001000",	-- 0x208b
		"00000101",	-- 0x208c
		"01010011",	-- 0x208d
		"00110111",	-- 0x208e
		"00010110",	-- 0x208f
		"00000001",	-- 0x2090
		"01010001",	-- 0x2091
		"01110101",	-- 0x2092
		"00011101",	-- 0x2093
		"00110011",	-- 0x2094
		"11111111",	-- 0x2095
		"10101001",	-- 0x2096
		"01110010",	-- 0x2097
		"10101000",	-- 0x2098
		"10110011",	-- 0x2099
		"00000001",	-- 0x209a
		"10000011",	-- 0x209b
		"01001010",	-- 0x209c
		"00000011",	-- 0x209d
		"01110101",	-- 0x209e
		"00101001",	-- 0x209f
		"10001100",	-- 0x20a0
		"01110111",	-- 0x20a1
		"00101001",	-- 0x20a2
		"01000000",	-- 0x20a3
		"01101100",	-- 0x20a4
		"10001111",	-- 0x20a5
		"11100000",	-- 0x20a6
		"11001100",	-- 0x20a7
		"11000000",	-- 0x20a8
		"00000011",	-- 0x20a9
		"00001101",	-- 0x20aa
		"11001100",	-- 0x20ab
		"01000010",	-- 0x20ac
		"01000010",	-- 0x20ad
		"00011101",	-- 0x20ae
		"10001110",	-- 0x20af
		"00000000",	-- 0x20b0
		"00000000",	-- 0x20b1
		"11101011",	-- 0x20b2
		"10000000",	-- 0x20b3
		"00001110",	-- 0x20b4
		"11101011",	-- 0x20b5
		"10000001",	-- 0x20b6
		"11101111",	-- 0x20b7
		"00000000",	-- 0x20b8
		"01000111",	-- 0x20b9
		"11101010",	-- 0x20ba
		"11001100",	-- 0x20bb
		"01000010",	-- 0x20bc
		"01000100",	-- 0x20bd
		"00001110",	-- 0x20be
		"11101011",	-- 0x20bf
		"10000010",	-- 0x20c0
		"11101101",	-- 0x20c1
		"10000101",	-- 0x20c2
		"01000110",	-- 0x20c3
		"00001000",	-- 0x20c4
		"11000000",	-- 0x20c5
		"00000011",	-- 0x20c6
		"00011101",	-- 0x20c7
		"00011101",	-- 0x20c8
		"00011101",	-- 0x20c9
		"01000000",	-- 0x20ca
		"11101111",	-- 0x20cb
		"01010010",	-- 0x20cc
		"01011000",	-- 0x20cd
		"01100011",	-- 0x20ce
		"10000000",	-- 0x20cf
		"00000001",	-- 0x20d0
		"00100001",	-- 0x20d1
		"10000000",	-- 0x20d2
		"10000000",	-- 0x20d3
		"00100001",	-- 0x20d4
		"10000000",	-- 0x20d5
		"00000010",	-- 0x20d6
		"00110001",	-- 0x20d7
		"10000000",	-- 0x20d8
		"00000100",	-- 0x20d9
		"01000001",	-- 0x20da
		"01101101",	-- 0x20db
		"00000001",	-- 0x20dc
		"01100001",	-- 0x20dd
		"10000010",	-- 0x20de
		"00100000",	-- 0x20df
		"00010010",	-- 0x20e0
		"10000010",	-- 0x20e1
		"00000100",	-- 0x20e2
		"00010010",	-- 0x20e3
		"10000000",	-- 0x20e4
		"00001000",	-- 0x20e5
		"00100010",	-- 0x20e6
		"10000010",	-- 0x20e7
		"00010000",	-- 0x20e8
		"00110010",	-- 0x20e9
		"10000000",	-- 0x20ea
		"00010000",	-- 0x20eb
		"01000010",	-- 0x20ec
		"10000010",	-- 0x20ed
		"01000000",	-- 0x20ee
		"01010010",	-- 0x20ef
		"10000000",	-- 0x20f0
		"00100000",	-- 0x20f1
		"00010011",	-- 0x20f2
		"10000100",	-- 0x20f3
		"00000001",	-- 0x20f4
		"01000011",	-- 0x20f5
		"10000010",	-- 0x20f6
		"00000010",	-- 0x20f7
		"00010100",	-- 0x20f8
		"10000000",	-- 0x20f9
		"01000000",	-- 0x20fa
		"00100100",	-- 0x20fb
		"10100000",	-- 0x20fc
		"00000100",	-- 0x20fd
		"00100100",	-- 0x20fe
		"10100000",	-- 0x20ff
		"00001000",	-- 0x2100
		"00110100",	-- 0x2101
		"10000010",	-- 0x2102
		"00001000",	-- 0x2103
		"01110100",	-- 0x2104
		"01001000",	-- 0x2105
		"00100000",	-- 0x2106
		"00010101",	-- 0x2107
		"10000010",	-- 0x2108
		"00000001",	-- 0x2109
		"00100101",	-- 0x210a
		"01001000",	-- 0x210b
		"00010000",	-- 0x210c
		"00110101",	-- 0x210d
		"10000010",	-- 0x210e
		"10000000",	-- 0x210f
		"01000101",	-- 0x2110
		"01100011",	-- 0x2111
		"00000011",	-- 0x2112
		"11100011",	-- 0x2113
		"01100011",	-- 0x2114
		"00110111",	-- 0x2115
		"10111001",	-- 0x2116
		"00100101",	-- 0x2117
		"00110111",	-- 0x2118
		"00011001",	-- 0x2119
		"00100100",	-- 0x211a
		"00110111",	-- 0x211b
		"01111001",	-- 0x211c
		"00100001",	-- 0x211d
		"00110111",	-- 0x211e
		"01011001",	-- 0x211f
		"00011110",	-- 0x2120
		"11111010",	-- 0x2121
		"00000001",	-- 0x2122
		"01010100",	-- 0x2123
		"11001100",	-- 0x2124
		"10011010",	-- 0x2125
		"01000101",	-- 0x2126
		"00010111",	-- 0x2127
		"11111010",	-- 0x2128
		"00000001",	-- 0x2129
		"01001111",	-- 0x212a
		"11001100",	-- 0x212b
		"10011010",	-- 0x212c
		"01000101",	-- 0x212d
		"00010000",	-- 0x212e
		"10010110",	-- 0x212f
		"01011001",	-- 0x2130
		"01000110",	-- 0x2131
		"00001100",	-- 0x2132
		"01111001",	-- 0x2133
		"10110100",	-- 0x2134
		"01011101",	-- 0x2135
		"01000101",	-- 0x2136
		"00000111",	-- 0x2137
		"00110101",	-- 0x2138
		"00111001",	-- 0x2139
		"00000111",	-- 0x213a
		"01000000",	-- 0x213b
		"00000010",	-- 0x213c
		"01110101",	-- 0x213d
		"00010000",	-- 0x213e
		"00000011",	-- 0x213f
		"11100010",	-- 0x2140
		"10110101",	-- 0x2141
		"01010010",	-- 0x2142
		"11001011",	-- 0x2143
		"00000100",	-- 0x2144
		"10011010",	-- 0x2145
		"00101110",	-- 0x2146
		"01110010",	-- 0x2147
		"00100111",	-- 0x2148
		"00110101",	-- 0x2149
		"11111001",	-- 0x214a
		"00011010",	-- 0x214b
		"00110101",	-- 0x214c
		"10011001",	-- 0x214d
		"00000011",	-- 0x214e
		"00000011",	-- 0x214f
		"11100001",	-- 0x2150
		"10011101",	-- 0x2151
		"11001010",	-- 0x2152
		"00001010",	-- 0x2153
		"10110010",	-- 0x2154
		"00000010",	-- 0x2155
		"00100011",	-- 0x2156
		"11001011",	-- 0x2157
		"00010101",	-- 0x2158
		"11000111",	-- 0x2159
		"11000000",	-- 0x215a
		"10110011",	-- 0x215b
		"00000010",	-- 0x215c
		"00100100",	-- 0x215d
		"00110011",	-- 0x215e
		"00000001",	-- 0x215f
		"00101001",	-- 0x2160
		"00110011",	-- 0x2161
		"00001101",	-- 0x2162
		"00100110",	-- 0x2163
		"01000000",	-- 0x2164
		"00100110",	-- 0x2165
		"11001010",	-- 0x2166
		"00010101",	-- 0x2167
		"00110111",	-- 0x2168
		"10101001",	-- 0x2169
		"00000010",	-- 0x216a
		"11001000",	-- 0x216b
		"00000001",	-- 0x216c
		"00110101",	-- 0x216d
		"11100010",	-- 0x216e
		"00000010",	-- 0x216f
		"11001000",	-- 0x2170
		"00000100",	-- 0x2171
		"10110010",	-- 0x2172
		"00000010",	-- 0x2173
		"00100011",	-- 0x2174
		"11001010",	-- 0x2175
		"00001010",	-- 0x2176
		"11000110",	-- 0x2177
		"10100000",	-- 0x2178
		"00110111",	-- 0x2179
		"00111010",	-- 0x217a
		"00000010",	-- 0x217b
		"11001000",	-- 0x217c
		"00000100",	-- 0x217d
		"00110111",	-- 0x217e
		"00011010",	-- 0x217f
		"00000010",	-- 0x2180
		"11001000",	-- 0x2181
		"00001000",	-- 0x2182
		"10110010",	-- 0x2183
		"00000010",	-- 0x2184
		"00100100",	-- 0x2185
		"00110011",	-- 0x2186
		"00000010",	-- 0x2187
		"00101001",	-- 0x2188
		"00110011",	-- 0x2189
		"00001110",	-- 0x218a
		"00100110",	-- 0x218b
		"10001110",	-- 0x218c
		"11111001",	-- 0x218d
		"11001000",	-- 0x218e
		"00011100",	-- 0x218f
		"01000110",	-- 0x2190
		"11111101",	-- 0x2191
		"00000001",	-- 0x2192
		"11100010",	-- 0x2193
		"01010100",	-- 0x2194
		"10001110",	-- 0x2195
		"11111001",	-- 0x2196
		"11000000",	-- 0x2197
		"00011100",	-- 0x2198
		"01000110",	-- 0x2199
		"11111101",	-- 0x219a
		"01000000",	-- 0x219b
		"10101100",	-- 0x219c
		"00000101",	-- 0x219d
		"01010010",	-- 0x219e
		"01010011",	-- 0x219f
		"10011010",	-- 0x21a0
		"00101110",	-- 0x21a1
		"11001010",	-- 0x21a2
		"10000000",	-- 0x21a3
		"10110010",	-- 0x21a4
		"00000010",	-- 0x21a5
		"00100100",	-- 0x21a6
		"10001110",	-- 0x21a7
		"11111001",	-- 0x21a8
		"11001000",	-- 0x21a9
		"00011100",	-- 0x21aa
		"01000110",	-- 0x21ab
		"11111101",	-- 0x21ac
		"00000001",	-- 0x21ad
		"11100010",	-- 0x21ae
		"01010100",	-- 0x21af
		"10001110",	-- 0x21b0
		"11111001",	-- 0x21b1
		"11000000",	-- 0x21b2
		"00011100",	-- 0x21b3
		"01000110",	-- 0x21b4
		"11111101",	-- 0x21b5
		"00000001",	-- 0x21b6
		"11100010",	-- 0x21b7
		"01101111",	-- 0x21b8
		"10001110",	-- 0x21b9
		"11111001",	-- 0x21ba
		"11000000",	-- 0x21bb
		"00011100",	-- 0x21bc
		"01000110",	-- 0x21bd
		"11111101",	-- 0x21be
		"00110011",	-- 0x21bf
		"00000100",	-- 0x21c0
		"00100010",	-- 0x21c1
		"00110011",	-- 0x21c2
		"00001000",	-- 0x21c3
		"00100110",	-- 0x21c4
		"10000101",	-- 0x21c5
		"00000000",	-- 0x21c6
		"10000101",	-- 0x21c7
		"00000000",	-- 0x21c8
		"01110101",	-- 0x21c9
		"01000111",	-- 0x21ca
		"01110111",	-- 0x21cb
		"01000110",	-- 0x21cc
		"11001011",	-- 0x21cd
		"00101111",	-- 0x21ce
		"01010001",	-- 0x21cf
		"01000110",	-- 0x21d0
		"11111101",	-- 0x21d1
		"01010111",	-- 0x21d2
		"00110011",	-- 0x21d3
		"00000011",	-- 0x21d4
		"00100010",	-- 0x21d5
		"00110111",	-- 0x21d6
		"10100010",	-- 0x21d7
		"00000110",	-- 0x21d8
		"00110101",	-- 0x21d9
		"10000010",	-- 0x21da
		"00000011",	-- 0x21db
		"00110101",	-- 0x21dc
		"01100010",	-- 0x21dd
		"00000010",	-- 0x21de
		"01000000",	-- 0x21df
		"01001111",	-- 0x21e0
		"01110101",	-- 0x21e1
		"00101001",	-- 0x21e2
		"01010010",	-- 0x21e3
		"01011011",	-- 0x21e4
		"10001111",	-- 0x21e5
		"00000000",	-- 0x21e6
		"01000000",	-- 0x21e7
		"10000010",	-- 0x21e8
		"01010110",	-- 0x21e9
		"10001101",	-- 0x21ea
		"00000011",	-- 0x21eb
		"00000000",	-- 0x21ec
		"01000101",	-- 0x21ed
		"11111001",	-- 0x21ee
		"10001111",	-- 0x21ef
		"00000000",	-- 0x21f0
		"01000000",	-- 0x21f1
		"00011010",	-- 0x21f2
		"00001011",	-- 0x21f3
		"01000110",	-- 0x21f4
		"00111001",	-- 0x21f5
		"01010111",	-- 0x21f6
		"10001101",	-- 0x21f7
		"00000011",	-- 0x21f8
		"00000000",	-- 0x21f9
		"01000101",	-- 0x21fa
		"11110110",	-- 0x21fb
		"00000001",	-- 0x21fc
		"11100010",	-- 0x21fd
		"01101111",	-- 0x21fe
		"01010111",	-- 0x21ff
		"01011010",	-- 0x2200
		"01000110",	-- 0x2201
		"11100001",	-- 0x2202
		"10001110",	-- 0x2203
		"11000000",	-- 0x2204
		"00000000",	-- 0x2205
		"01010010",	-- 0x2206
		"01010011",	-- 0x2207
		"10001111",	-- 0x2208
		"00000001",	-- 0x2209
		"00000000",	-- 0x220a
		"10100111",	-- 0x220b
		"00000000",	-- 0x220c
		"00011100",	-- 0x220d
		"00011100",	-- 0x220e
		"00011111",	-- 0x220f
		"01000110",	-- 0x2210
		"11111001",	-- 0x2211
		"00000001",	-- 0x2212
		"11100010",	-- 0x2213
		"01101111",	-- 0x2214
		"10001100",	-- 0x2215
		"00000000",	-- 0x2216
		"00000000",	-- 0x2217
		"01000110",	-- 0x2218
		"11101110",	-- 0x2219
		"10001001",	-- 0x221a
		"10101010",	-- 0x221b
		"01010101",	-- 0x221c
		"01000110",	-- 0x221d
		"00010000",	-- 0x221e
		"00110101",	-- 0x221f
		"10100010",	-- 0x2220
		"00001110",	-- 0x2221
		"00110111",	-- 0x2222
		"10000010",	-- 0x2223
		"00001011",	-- 0x2224
		"00110101",	-- 0x2225
		"01100010",	-- 0x2226
		"00001000",	-- 0x2227
		"00010011",	-- 0x2228
		"01110111",	-- 0x2229
		"00101001",	-- 0x222a
		"11001010",	-- 0x222b
		"00011001",	-- 0x222c
		"01000000",	-- 0x222d
		"00010011",	-- 0x222e
		"01010011",	-- 0x222f
		"01110001",	-- 0x2230
		"00101001",	-- 0x2231
		"01000111",	-- 0x2232
		"00000010",	-- 0x2233
		"01110101",	-- 0x2234
		"00101001",	-- 0x2235
		"11001010",	-- 0x2236
		"01111101",	-- 0x2237
		"01011001",	-- 0x2238
		"01000111",	-- 0x2239
		"00000111",	-- 0x223a
		"11001101",	-- 0x223b
		"11111111",	-- 0x223c
		"01000110",	-- 0x223d
		"00000010",	-- 0x223e
		"11001010",	-- 0x223f
		"01011110",	-- 0x2240
		"00010010",	-- 0x2241
		"10001110",	-- 0x2242
		"11110111",	-- 0x2243
		"10110101",	-- 0x2244
		"00011100",	-- 0x2245
		"01000110",	-- 0x2246
		"11111101",	-- 0x2247
		"01100001",	-- 0x2248
		"00100101",	-- 0x2249
		"01010000",	-- 0x224a
		"01000110",	-- 0x224b
		"11110101",	-- 0x224c
		"11001101",	-- 0x224d
		"10101010",	-- 0x224e
		"01000110",	-- 0x224f
		"11011111",	-- 0x2250
		"00000011",	-- 0x2251
		"11100001",	-- 0x2252
		"11100001",	-- 0x2253
		"01101000",	-- 0x2254
		"01110001",	-- 0x2255
		"00000000",	-- 0x2256
		"01000111",	-- 0x2257
		"00000010",	-- 0x2258
		"01110101",	-- 0x2259
		"00000000",	-- 0x225a
		"00000001",	-- 0x225b
		"11111011",	-- 0x225c
		"00011101",	-- 0x225d
		"00000001",	-- 0x225e
		"11111000",	-- 0x225f
		"01111100",	-- 0x2260
		"00110111",	-- 0x2261
		"00011001",	-- 0x2262
		"00011110",	-- 0x2263
		"00110111",	-- 0x2264
		"01111001",	-- 0x2265
		"00011011",	-- 0x2266
		"00110101",	-- 0x2267
		"11000010",	-- 0x2268
		"00011000",	-- 0x2269
		"00110101",	-- 0x226a
		"01000000",	-- 0x226b
		"00010101",	-- 0x226c
		"01111000",	-- 0x226d
		"01100011",	-- 0x226e
		"01110001",	-- 0x226f
		"00000000",	-- 0x2270
		"01000111",	-- 0x2271
		"00000010",	-- 0x2272
		"01110101",	-- 0x2273
		"00000000",	-- 0x2274
		"00110111",	-- 0x2275
		"00100000",	-- 0x2276
		"00001010",	-- 0x2277
		"00110101",	-- 0x2278
		"10000000",	-- 0x2279
		"00000111",	-- 0x227a
		"00110101",	-- 0x227b
		"11000010",	-- 0x227c
		"00000100",	-- 0x227d
		"00110101",	-- 0x227e
		"01000000",	-- 0x227f
		"00000001",	-- 0x2280
		"01100011",	-- 0x2281
		"10001110",	-- 0x2282
		"11111001",	-- 0x2283
		"11000000",	-- 0x2284
		"00011100",	-- 0x2285
		"01000110",	-- 0x2286
		"11111101",	-- 0x2287
		"01110001",	-- 0x2288
		"00000000",	-- 0x2289
		"01000111",	-- 0x228a
		"00000010",	-- 0x228b
		"01110101",	-- 0x228c
		"00000000",	-- 0x228d
		"10001110",	-- 0x228e
		"11111001",	-- 0x228f
		"11000000",	-- 0x2290
		"00011100",	-- 0x2291
		"01000110",	-- 0x2292
		"11111101",	-- 0x2293
		"10001111",	-- 0x2294
		"00000000",	-- 0x2295
		"01000000",	-- 0x2296
		"01010010",	-- 0x2297
		"01010011",	-- 0x2298
		"10011010",	-- 0x2299
		"00101100",	-- 0x229a
		"10001010",	-- 0x229b
		"10001101",	-- 0x229c
		"00000010",	-- 0x229d
		"11111111",	-- 0x229e
		"01000011",	-- 0x229f
		"11111010",	-- 0x22a0
		"10001011",	-- 0x22a1
		"00000010",	-- 0x22a2
		"11111111",	-- 0x22a3
		"00110011",	-- 0x22a4
		"11011101",	-- 0x22a5
		"00100000",	-- 0x22a6
		"00110011",	-- 0x22a7
		"11011001",	-- 0x22a8
		"00100010",	-- 0x22a9
		"00110011",	-- 0x22aa
		"00000011",	-- 0x22ab
		"00101001",	-- 0x22ac
		"00110011",	-- 0x22ad
		"00001000",	-- 0x22ae
		"00100110",	-- 0x22af
		"01110111",	-- 0x22b0
		"00010000",	-- 0x22b1
		"00000011",	-- 0x22b2
		"11000110",	-- 0x22b3
		"01111010",	-- 0x22b4
		"00110101",	-- 0x22b5
		"00010000",	-- 0x22b6
		"00000011",	-- 0x22b7
		"00000011",	-- 0x22b8
		"11100011",	-- 0x22b9
		"01100010",	-- 0x22ba
		"11001010",	-- 0x22bb
		"00001001",	-- 0x22bc
		"11000110",	-- 0x22bd
		"11100000",	-- 0x22be
		"10110010",	-- 0x22bf
		"00000010",	-- 0x22c0
		"00100100",	-- 0x22c1
		"01010010",	-- 0x22c2
		"00110101",	-- 0x22c3
		"00111001",	-- 0x22c4
		"00010110",	-- 0x22c5
		"00110111",	-- 0x22c6
		"11011010",	-- 0x22c7
		"00000010",	-- 0x22c8
		"11000110",	-- 0x22c9
		"00000001",	-- 0x22ca
		"00110111",	-- 0x22cb
		"11111010",	-- 0x22cc
		"00000010",	-- 0x22cd
		"11000110",	-- 0x22ce
		"00000010",	-- 0x22cf
		"00110111",	-- 0x22d0
		"01111010",	-- 0x22d1
		"00000010",	-- 0x22d2
		"11000110",	-- 0x22d3
		"00000100",	-- 0x22d4
		"00110111",	-- 0x22d5
		"01011010",	-- 0x22d6
		"00000010",	-- 0x22d7
		"11000110",	-- 0x22d8
		"00001000",	-- 0x22d9
		"01000000",	-- 0x22da
		"00010111",	-- 0x22db
		"00110111",	-- 0x22dc
		"10011010",	-- 0x22dd
		"00000010",	-- 0x22de
		"11000110",	-- 0x22df
		"00000001",	-- 0x22e0
		"00110111",	-- 0x22e1
		"10111010",	-- 0x22e2
		"00000010",	-- 0x22e3
		"11000110",	-- 0x22e4
		"00000010",	-- 0x22e5
		"00110111",	-- 0x22e6
		"01011001",	-- 0x22e7
		"00000010",	-- 0x22e8
		"11000110",	-- 0x22e9
		"00000100",	-- 0x22ea
		"11011011",	-- 0x22eb
		"00000111",	-- 0x22ec
		"11001111",	-- 0x22ed
		"00000010",	-- 0x22ee
		"01000111",	-- 0x22ef
		"00000010",	-- 0x22f0
		"11000110",	-- 0x22f1
		"00001000",	-- 0x22f2
		"11011011",	-- 0x22f3
		"01010111",	-- 0x22f4
		"11001101",	-- 0x22f5
		"00011000",	-- 0x22f6
		"01000101",	-- 0x22f7
		"01011111",	-- 0x22f8
		"11111010",	-- 0x22f9
		"00000010",	-- 0x22fa
		"01000101",	-- 0x22fb
		"11001101",	-- 0x22fc
		"00100110",	-- 0x22fd
		"01000101",	-- 0x22fe
		"01011101",	-- 0x22ff
		"11111010",	-- 0x2300
		"00000010",	-- 0x2301
		"01000100",	-- 0x2302
		"11001101",	-- 0x2303
		"00111010",	-- 0x2304
		"01000101",	-- 0x2305
		"01010011",	-- 0x2306
		"11111010",	-- 0x2307
		"00000001",	-- 0x2308
		"11001110",	-- 0x2309
		"00110111",	-- 0x230a
		"00011001",	-- 0x230b
		"00001111",	-- 0x230c
		"11111010",	-- 0x230d
		"00000001",	-- 0x230e
		"11001101",	-- 0x230f
		"00110111",	-- 0x2310
		"00111001",	-- 0x2311
		"00001001",	-- 0x2312
		"11111010",	-- 0x2313
		"00000001",	-- 0x2314
		"11001100",	-- 0x2315
		"00110111",	-- 0x2316
		"01111001",	-- 0x2317
		"00000011",	-- 0x2318
		"11111010",	-- 0x2319
		"00000001",	-- 0x231a
		"11001011",	-- 0x231b
		"11001101",	-- 0x231c
		"01101011",	-- 0x231d
		"01000101",	-- 0x231e
		"00111101",	-- 0x231f
		"11011010",	-- 0x2320
		"01010100",	-- 0x2321
		"00110111",	-- 0x2322
		"00111001",	-- 0x2323
		"00000011",	-- 0x2324
		"11111010",	-- 0x2325
		"00000010",	-- 0x2326
		"00101110",	-- 0x2327
		"11001101",	-- 0x2328
		"10010010",	-- 0x2329
		"01000101",	-- 0x232a
		"00110001",	-- 0x232b
		"11111010",	-- 0x232c
		"00000001",	-- 0x232d
		"01001111",	-- 0x232e
		"11001101",	-- 0x232f
		"10101001",	-- 0x2330
		"01000101",	-- 0x2331
		"00101010",	-- 0x2332
		"11111010",	-- 0x2333
		"00000001",	-- 0x2334
		"10000110",	-- 0x2335
		"11001101",	-- 0x2336
		"10111100",	-- 0x2337
		"01000101",	-- 0x2338
		"00100011",	-- 0x2339
		"11001010",	-- 0x233a
		"10111000",	-- 0x233b
		"11001101",	-- 0x233c
		"11001011",	-- 0x233d
		"01000101",	-- 0x233e
		"00011101",	-- 0x233f
		"11011010",	-- 0x2340
		"01011101",	-- 0x2341
		"11001101",	-- 0x2342
		"11011100",	-- 0x2343
		"01000101",	-- 0x2344
		"00010111",	-- 0x2345
		"11111010",	-- 0x2346
		"00000001",	-- 0x2347
		"00000010",	-- 0x2348
		"11001101",	-- 0x2349
		"11101010",	-- 0x234a
		"01000101",	-- 0x234b
		"00010000",	-- 0x234c
		"11011010",	-- 0x234d
		"01010101",	-- 0x234e
		"11001101",	-- 0x234f
		"11110011",	-- 0x2350
		"01000101",	-- 0x2351
		"00001010",	-- 0x2352
		"11111010",	-- 0x2353
		"00000001",	-- 0x2354
		"01010100",	-- 0x2355
		"01000000",	-- 0x2356
		"00000101",	-- 0x2357
		"11000000",	-- 0x2358
		"00001000",	-- 0x2359
		"00010010",	-- 0x235a
		"00010010",	-- 0x235b
		"00010010",	-- 0x235c
		"10000001",	-- 0x235d
		"00000100",	-- 0x235e
		"10111010",	-- 0x235f
		"00000001",	-- 0x2360
		"10011000",	-- 0x2361
		"01100011",	-- 0x2362
		"01110001",	-- 0x2363
		"11110001",	-- 0x2364
		"01000111",	-- 0x2365
		"00000011",	-- 0x2366
		"00000011",	-- 0x2367
		"11100011",	-- 0x2368
		"10100110",	-- 0x2369
		"10000110",	-- 0x236a
		"11100001",	-- 0x236b
		"00000111",	-- 0x236c
		"00000001",	-- 0x236d
		"11000100",	-- 0x236e
		"10111001",	-- 0x236f
		"11011010",	-- 0x2370
		"11101000",	-- 0x2371
		"01010110",	-- 0x2372
		"10010010",	-- 0x2373
		"11101000",	-- 0x2374
		"11001110",	-- 0x2375
		"00000001",	-- 0x2376
		"01000110",	-- 0x2377
		"00000110",	-- 0x2378
		"10000110",	-- 0x2379
		"11101001",	-- 0x237a
		"00000001",	-- 0x237b
		"00000001",	-- 0x237c
		"11000100",	-- 0x237d
		"10111001",	-- 0x237e
		"00000001",	-- 0x237f
		"11100100",	-- 0x2380
		"00110101",	-- 0x2381
		"00000001",	-- 0x2382
		"11001011",	-- 0x2383
		"00001011",	-- 0x2384
		"00000001",	-- 0x2385
		"11101100",	-- 0x2386
		"00011010",	-- 0x2387
		"00000001",	-- 0x2388
		"11010011",	-- 0x2389
		"01110110",	-- 0x238a
		"11111010",	-- 0x238b
		"00000001",	-- 0x238c
		"11010111",	-- 0x238d
		"10010010",	-- 0x238e
		"01001110",	-- 0x238f
		"00000001",	-- 0x2390
		"11010100",	-- 0x2391
		"10111100",	-- 0x2392
		"11111010",	-- 0x2393
		"00000001",	-- 0x2394
		"11010001",	-- 0x2395
		"10010010",	-- 0x2396
		"01001110",	-- 0x2397
		"00000001",	-- 0x2398
		"11011010",	-- 0x2399
		"01100011",	-- 0x239a
		"11011010",	-- 0x239b
		"01001110",	-- 0x239c
		"10110010",	-- 0x239d
		"00000001",	-- 0x239e
		"11010001",	-- 0x239f
		"00000001",	-- 0x23a0
		"11011101",	-- 0x23a1
		"01101001",	-- 0x23a2
		"00000001",	-- 0x23a3
		"11100001",	-- 0x23a4
		"00010101",	-- 0x23a5
		"00000001",	-- 0x23a6
		"11100100",	-- 0x23a7
		"01010100",	-- 0x23a8
		"00000001",	-- 0x23a9
		"11100101",	-- 0x23aa
		"01010001",	-- 0x23ab
		"00110101",	-- 0x23ac
		"00010110",	-- 0x23ad
		"00000011",	-- 0x23ae
		"00000011",	-- 0x23af
		"11100100",	-- 0x23b0
		"01010010",	-- 0x23b1
		"10001111",	-- 0x23b2
		"11000001",	-- 0x23b3
		"00010010",	-- 0x23b4
		"00000001",	-- 0x23b5
		"11000011",	-- 0x23b6
		"11101110",	-- 0x23b7
		"10011010",	-- 0x23b8
		"01111010",	-- 0x23b9
		"10010110",	-- 0x23ba
		"01011001",	-- 0x23bb
		"10001111",	-- 0x23bc
		"11000001",	-- 0x23bd
		"00101101",	-- 0x23be
		"00000001",	-- 0x23bf
		"11000100",	-- 0x23c0
		"00110100",	-- 0x23c1
		"01101100",	-- 0x23c2
		"10001111",	-- 0x23c3
		"11000001",	-- 0x23c4
		"00110111",	-- 0x23c5
		"00000001",	-- 0x23c6
		"11000100",	-- 0x23c7
		"01000010",	-- 0x23c8
		"01111101",	-- 0x23c9
		"00001011",	-- 0x23ca
		"01000100",	-- 0x23cb
		"00000001",	-- 0x23cc
		"01011011",	-- 0x23cd
		"00110101",	-- 0x23ce
		"00010000",	-- 0x23cf
		"00001000",	-- 0x23d0
		"11011010",	-- 0x23d1
		"10011111",	-- 0x23d2
		"11001100",	-- 0x23d3
		"01111010",	-- 0x23d4
		"01000101",	-- 0x23d5
		"00000010",	-- 0x23d6
		"11001011",	-- 0x23d7
		"00011010",	-- 0x23d8
		"01010010",	-- 0x23d9
		"10011110",	-- 0x23da
		"01111010",	-- 0x23db
		"00000001",	-- 0x23dc
		"11000101",	-- 0x23dd
		"00000111",	-- 0x23de
		"10011010",	-- 0x23df
		"01111010",	-- 0x23e0
		"11011011",	-- 0x23e1
		"01010110",	-- 0x23e2
		"10001111",	-- 0x23e3
		"11000001",	-- 0x23e4
		"00111100",	-- 0x23e5
		"00000001",	-- 0x23e6
		"11000100",	-- 0x23e7
		"01000111",	-- 0x23e8
		"01011011",	-- 0x23e9
		"10011110",	-- 0x23ea
		"01111010",	-- 0x23eb
		"00000001",	-- 0x23ec
		"11000101",	-- 0x23ed
		"01001111",	-- 0x23ee
		"10011010",	-- 0x23ef
		"01111010",	-- 0x23f0
		"00110111",	-- 0x23f1
		"11110110",	-- 0x23f2
		"00010001",	-- 0x23f3
		"10000110",	-- 0x23f4
		"00000111",	-- 0x23f5
		"01011000",	-- 0x23f6
		"00110101",	-- 0x23f7
		"00011001",	-- 0x23f8
		"00101001",	-- 0x23f9
		"10000110",	-- 0x23fa
		"00000101",	-- 0x23fb
		"01100100",	-- 0x23fc
		"00110111",	-- 0x23fd
		"01010110",	-- 0x23fe
		"00100011",	-- 0x23ff
		"10000110",	-- 0x2400
		"00000001",	-- 0x2401
		"01001010",	-- 0x2402
		"01000000",	-- 0x2403
		"00011110",	-- 0x2404
		"00110101",	-- 0x2405
		"01111101",	-- 0x2406
		"00010011",	-- 0x2407
		"01010011",	-- 0x2408
		"11011010",	-- 0x2409
		"10011000",	-- 0x240a
		"00110101",	-- 0x240b
		"00010010",	-- 0x240c
		"00000010",	-- 0x240d
		"11001010",	-- 0x240e
		"01010000",	-- 0x240f
		"10000101",	-- 0x2410
		"01100001",	-- 0x2411
		"01000100",	-- 0x2412
		"00000010",	-- 0x2413
		"11001011",	-- 0x2414
		"11111111",	-- 0x2415
		"10011110",	-- 0x2416
		"01111010",	-- 0x2417
		"00000001",	-- 0x2418
		"11000101",	-- 0x2419
		"01011010",	-- 0x241a
		"10001001",	-- 0x241b
		"11110100",	-- 0x241c
		"00100100",	-- 0x241d
		"01000011",	-- 0x241e
		"00000011",	-- 0x241f
		"10000110",	-- 0x2420
		"11110100",	-- 0x2421
		"00100100",	-- 0x2422
		"00000101",	-- 0x2423
		"10111010",	-- 0x2424
		"00000001",	-- 0x2425
		"00001010",	-- 0x2426
		"10111010",	-- 0x2427
		"00000001",	-- 0x2428
		"00001100",	-- 0x2429
		"10111010",	-- 0x242a
		"00000001",	-- 0x242b
		"00001110",	-- 0x242c
		"10111010",	-- 0x242d
		"00000001",	-- 0x242e
		"00010000",	-- 0x242f
		"01110101",	-- 0x2430
		"11110101",	-- 0x2431
		"00000111",	-- 0x2432
		"01000000",	-- 0x2433
		"00011101",	-- 0x2434
		"11011010",	-- 0x2435
		"10011111",	-- 0x2436
		"00110111",	-- 0x2437
		"00010110",	-- 0x2438
		"00000110",	-- 0x2439
		"00110111",	-- 0x243a
		"00011001",	-- 0x243b
		"00000011",	-- 0x243c
		"01010110",	-- 0x243d
		"01000111",	-- 0x243e
		"00001110",	-- 0x243f
		"01111001",	-- 0x2440
		"00100000",	-- 0x2441
		"01011011",	-- 0x2442
		"01000100",	-- 0x2443
		"00001001",	-- 0x2444
		"01111001",	-- 0x2445
		"00111101",	-- 0x2446
		"11010000",	-- 0x2447
		"01000100",	-- 0x2448
		"00000100",	-- 0x2449
		"11001100",	-- 0x244a
		"10101000",	-- 0x244b
		"01000101",	-- 0x244c
		"00000001",	-- 0x244d
		"01010010",	-- 0x244e
		"10010010",	-- 0x244f
		"10011111",	-- 0x2450
		"01100011",	-- 0x2451
		"01000000",	-- 0x2452
		"01100101",	-- 0x2453
		"10111110",	-- 0x2454
		"00000001",	-- 0x2455
		"00111010",	-- 0x2456
		"11111010",	-- 0x2457
		"00000010",	-- 0x2458
		"00110111",	-- 0x2459
		"01000111",	-- 0x245a
		"00010111",	-- 0x245b
		"00110111",	-- 0x245c
		"01010100",	-- 0x245d
		"00001010",	-- 0x245e
		"00110111",	-- 0x245f
		"01011101",	-- 0x2460
		"00000111",	-- 0x2461
		"10000001",	-- 0x2462
		"10000000",	-- 0x2463
		"00000110",	-- 0x2464
		"01000100",	-- 0x2465
		"00000010",	-- 0x2466
		"11001010",	-- 0x2467
		"11111111",	-- 0x2468
		"01011011",	-- 0x2469
		"11000001",	-- 0x246a
		"10000000",	-- 0x246b
		"01000100",	-- 0x246c
		"00000010",	-- 0x246d
		"11001011",	-- 0x246e
		"11111111",	-- 0x246f
		"00000001",	-- 0x2470
		"11000101",	-- 0x2471
		"01001111",	-- 0x2472
		"11111011",	-- 0x2473
		"00000001",	-- 0x2474
		"00011100",	-- 0x2475
		"01001011",	-- 0x2476
		"00000011",	-- 0x2477
		"00000001",	-- 0x2478
		"11000101",	-- 0x2479
		"01001111",	-- 0x247a
		"01101110",	-- 0x247b
		"00000001",	-- 0x247c
		"11010001",	-- 0x247d
		"10100001",	-- 0x247e
		"01010010",	-- 0x247f
		"11010001",	-- 0x2480
		"01100010",	-- 0x2481
		"10000000",	-- 0x2482
		"00000000",	-- 0x2483
		"10000111",	-- 0x2484
		"00000001",	-- 0x2485
		"00000000",	-- 0x2486
		"10011010",	-- 0x2487
		"01111000",	-- 0x2488
		"00101110",	-- 0x2489
		"10101110",	-- 0x248a
		"00000000",	-- 0x248b
		"00000001",	-- 0x248c
		"11000100",	-- 0x248d
		"11110101",	-- 0x248e
		"00000001",	-- 0x248f
		"11000100",	-- 0x2490
		"11011100",	-- 0x2491
		"10110011",	-- 0x2492
		"00000001",	-- 0x2493
		"11001010",	-- 0x2494
		"11111010",	-- 0x2495
		"00000001",	-- 0x2496
		"11010001",	-- 0x2497
		"10010010",	-- 0x2498
		"01001110",	-- 0x2499
		"00000001",	-- 0x249a
		"11011011",	-- 0x249b
		"10100011",	-- 0x249c
		"11011010",	-- 0x249d
		"01001110",	-- 0x249e
		"10110010",	-- 0x249f
		"00000001",	-- 0x24a0
		"11010001",	-- 0x24a1
		"10110110",	-- 0x24a2
		"00000001",	-- 0x24a3
		"11000110",	-- 0x24a4
		"00000001",	-- 0x24a5
		"11000100",	-- 0x24a6
		"11001001",	-- 0x24a7
		"10010111",	-- 0x24a8
		"01111000",	-- 0x24a9
		"10001000",	-- 0x24aa
		"00000001",	-- 0x24ab
		"10011001",	-- 0x24ac
		"01000100",	-- 0x24ad
		"00000010",	-- 0x24ae
		"01010010",	-- 0x24af
		"01010011",	-- 0x24b0
		"01111110",	-- 0x24b1
		"00000001",	-- 0x24b2
		"11000100",	-- 0x24b3
		"11110101",	-- 0x24b4
		"10111010",	-- 0x24b5
		"00000001",	-- 0x24b6
		"00111000",	-- 0x24b7
		"01100011",	-- 0x24b8
		"10001110",	-- 0x24b9
		"00000000",	-- 0x24ba
		"10000000",	-- 0x24bb
		"11111010",	-- 0x24bc
		"00000010",	-- 0x24bd
		"00110000",	-- 0x24be
		"00001100",	-- 0x24bf
		"11111010",	-- 0x24c0
		"00000010",	-- 0x24c1
		"00110001",	-- 0x24c2
		"00001100",	-- 0x24c3
		"00001100",	-- 0x24c4
		"11111010",	-- 0x24c5
		"00000010",	-- 0x24c6
		"00110100",	-- 0x24c7
		"00001100",	-- 0x24c8
		"00001100",	-- 0x24c9
		"00001100",	-- 0x24ca
		"00001100",	-- 0x24cb
		"00110111",	-- 0x24cc
		"01010110",	-- 0x24cd
		"00000101",	-- 0x24ce
		"11111010",	-- 0x24cf
		"00000010",	-- 0x24d0
		"00110011",	-- 0x24d1
		"00001100",	-- 0x24d2
		"00001100",	-- 0x24d3
		"11111010",	-- 0x24d4
		"00000010",	-- 0x24d5
		"00110110",	-- 0x24d6
		"00001100",	-- 0x24d7
		"00111100",	-- 0x24d8
		"11110101",	-- 0x24d9
		"00000001",	-- 0x24da
		"00100000",	-- 0x24db
		"10000100",	-- 0x24dc
		"00000000",	-- 0x24dd
		"00000110",	-- 0x24de
		"00111110",	-- 0x24df
		"11111011",	-- 0x24e0
		"00000010",	-- 0x24e1
		"00111011",	-- 0x24e2
		"11001101",	-- 0x24e3
		"10000000",	-- 0x24e4
		"01000111",	-- 0x24e5
		"00000100",	-- 0x24e6
		"00000001",	-- 0x24e7
		"11000100",	-- 0x24e8
		"11110001",	-- 0x24e9
		"00111110",	-- 0x24ea
		"10110110",	-- 0x24eb
		"00000010",	-- 0x24ec
		"00101100",	-- 0x24ed
		"00000001",	-- 0x24ee
		"11000101",	-- 0x24ef
		"00000111",	-- 0x24f0
		"00111110",	-- 0x24f1
		"00110111",	-- 0x24f2
		"01010110",	-- 0x24f3
		"00000101",	-- 0x24f4
		"11011011",	-- 0x24f5
		"01100000",	-- 0x24f6
		"00000001",	-- 0x24f7
		"11000101",	-- 0x24f8
		"01001111",	-- 0x24f9
		"11111011",	-- 0x24fa
		"00000010",	-- 0x24fb
		"00110101",	-- 0x24fc
		"00000001",	-- 0x24fd
		"11000100",	-- 0x24fe
		"11110001",	-- 0x24ff
		"10111010",	-- 0x2500
		"00000001",	-- 0x2501
		"00111010",	-- 0x2502
		"01110101",	-- 0x2503
		"00011000",	-- 0x2504
		"11011010",	-- 0x2505
		"10011010",	-- 0x2506
		"00110101",	-- 0x2507
		"00010010",	-- 0x2508
		"00000010",	-- 0x2509
		"11001010",	-- 0x250a
		"01100110",	-- 0x250b
		"10000001",	-- 0x250c
		"00000100",	-- 0x250d
		"10011010",	-- 0x250e
		"01111001",	-- 0x250f
		"10110110",	-- 0x2510
		"00000001",	-- 0x2511
		"10011000",	-- 0x2512
		"10011000",	-- 0x2513
		"01111001",	-- 0x2514
		"01000100",	-- 0x2515
		"00000011",	-- 0x2516
		"00000001",	-- 0x2517
		"11000100",	-- 0x2518
		"11100111",	-- 0x2519
		"00111110",	-- 0x251a
		"11001010",	-- 0x251b
		"00011001",	-- 0x251c
		"00000001",	-- 0x251d
		"11000101",	-- 0x251e
		"01011011",	-- 0x251f
		"00000001",	-- 0x2520
		"11000100",	-- 0x2521
		"11101001",	-- 0x2522
		"00110111",	-- 0x2523
		"00111000",	-- 0x2524
		"00000101",	-- 0x2525
		"10000111",	-- 0x2526
		"00000000",	-- 0x2527
		"00010000",	-- 0x2528
		"01001001",	-- 0x2529
		"00000101",	-- 0x252a
		"01011000",	-- 0x252b
		"01001011",	-- 0x252c
		"00000101",	-- 0x252d
		"01000111",	-- 0x252e
		"00000100",	-- 0x252f
		"11001011",	-- 0x2530
		"11111111",	-- 0x2531
		"01000001",	-- 0x2532
		"01010011",	-- 0x2533
		"10110011",	-- 0x2534
		"00000001",	-- 0x2535
		"01000011",	-- 0x2536
		"01000000",	-- 0x2537
		"00010101",	-- 0x2538
		"10010110",	-- 0x2539
		"01010010",	-- 0x253a
		"01011000",	-- 0x253b
		"01000110",	-- 0x253c
		"00000001",	-- 0x253d
		"01010011",	-- 0x253e
		"10011010",	-- 0x253f
		"01111000",	-- 0x2540
		"11111010",	-- 0x2541
		"00000001",	-- 0x2542
		"01000011",	-- 0x2543
		"10000001",	-- 0x2544
		"01000000",	-- 0x2545
		"10010111",	-- 0x2546
		"01111000",	-- 0x2547
		"01000100",	-- 0x2548
		"00000011",	-- 0x2549
		"10000110",	-- 0x254a
		"11111111",	-- 0x254b
		"11111111",	-- 0x254c
		"01100011",	-- 0x254d
		"00000011",	-- 0x254e
		"11100111",	-- 0x254f
		"11001101",	-- 0x2550
		"00000001",	-- 0x2551
		"11100111",	-- 0x2552
		"01100111",	-- 0x2553
		"10110010",	-- 0x2554
		"00000001",	-- 0x2555
		"00110111",	-- 0x2556
		"00111100",	-- 0x2557
		"10110010",	-- 0x2558
		"00000001",	-- 0x2559
		"01000101",	-- 0x255a
		"11111011",	-- 0x255b
		"00000001",	-- 0x255c
		"01000100",	-- 0x255d
		"00000001",	-- 0x255e
		"11000101",	-- 0x255f
		"01001111",	-- 0x2560
		"00001010",	-- 0x2561
		"00000001",	-- 0x2562
		"00110001",	-- 0x2563
		"10010110",	-- 0x2564
		"01010000",	-- 0x2565
		"00110101",	-- 0x2566
		"00010000",	-- 0x2567
		"00000110",	-- 0x2568
		"00110101",	-- 0x2569
		"00010110",	-- 0x256a
		"00000011",	-- 0x256b
		"00110111",	-- 0x256c
		"11110111",	-- 0x256d
		"00000011",	-- 0x256e
		"00000011",	-- 0x256f
		"11100110",	-- 0x2570
		"00100111",	-- 0x2571
		"10110110",	-- 0x2572
		"00000001",	-- 0x2573
		"00001010",	-- 0x2574
		"10000111",	-- 0x2575
		"00000101",	-- 0x2576
		"10010001",	-- 0x2577
		"01000100",	-- 0x2578
		"00000011",	-- 0x2579
		"10000110",	-- 0x257a
		"11111111",	-- 0x257b
		"11111111",	-- 0x257c
		"00000100",	-- 0x257d
		"00000100",	-- 0x257e
		"00000100",	-- 0x257f
		"10011010",	-- 0x2580
		"01111000",	-- 0x2581
		"11111010",	-- 0x2582
		"00000001",	-- 0x2583
		"00001001",	-- 0x2584
		"10000001",	-- 0x2585
		"10101011",	-- 0x2586
		"10000111",	-- 0x2587
		"00000101",	-- 0x2588
		"00111111",	-- 0x2589
		"01000100",	-- 0x258a
		"00000011",	-- 0x258b
		"10000110",	-- 0x258c
		"11111111",	-- 0x258d
		"11111111",	-- 0x258e
		"10001000",	-- 0x258f
		"00000111",	-- 0x2590
		"01010101",	-- 0x2591
		"00000001",	-- 0x2592
		"11000100",	-- 0x2593
		"11011100",	-- 0x2594
		"01011010",	-- 0x2595
		"10001111",	-- 0x2596
		"00000000",	-- 0x2597
		"11110110",	-- 0x2598
		"10100001",	-- 0x2599
		"10000000",	-- 0x259a
		"10000111",	-- 0x259b
		"00000001",	-- 0x259c
		"00000000",	-- 0x259d
		"01000101",	-- 0x259e
		"00000100",	-- 0x259f
		"10010111",	-- 0x25a0
		"01111000",	-- 0x25a1
		"01000100",	-- 0x25a2
		"00000010",	-- 0x25a3
		"11001010",	-- 0x25a4
		"11111111",	-- 0x25a5
		"11001100",	-- 0x25a6
		"00001110",	-- 0x25a7
		"01000011",	-- 0x25a8
		"00000010",	-- 0x25a9
		"11001010",	-- 0x25aa
		"00001110",	-- 0x25ab
		"01101100",	-- 0x25ac
		"00010000",	-- 0x25ad
		"10010010",	-- 0x25ae
		"01111011",	-- 0x25af
		"00110111",	-- 0x25b0
		"11010111",	-- 0x25b1
		"00101001",	-- 0x25b2
		"01100001",	-- 0x25b3
		"10000100",	-- 0x25b4
		"00000001",	-- 0x25b5
		"11000100",	-- 0x25b6
		"11001010",	-- 0x25b7
		"10011010",	-- 0x25b8
		"01111000",	-- 0x25b9
		"11011010",	-- 0x25ba
		"01011110",	-- 0x25bb
		"10010010",	-- 0x25bc
		"01111010",	-- 0x25bd
		"10010001",	-- 0x25be
		"01111011",	-- 0x25bf
		"01111001",	-- 0x25c0
		"00000000",	-- 0x25c1
		"01111010",	-- 0x25c2
		"01001010",	-- 0x25c3
		"00001001",	-- 0x25c4
		"11010100",	-- 0x25c5
		"01111011",	-- 0x25c6
		"10010111",	-- 0x25c7
		"01111000",	-- 0x25c8
		"01000101",	-- 0x25c9
		"00000101",	-- 0x25ca
		"01010010",	-- 0x25cb
		"01010011",	-- 0x25cc
		"10001100",	-- 0x25cd
		"10010111",	-- 0x25ce
		"01111000",	-- 0x25cf
		"00000110",	-- 0x25d0
		"00000110",	-- 0x25d1
		"00000110",	-- 0x25d2
		"00000001",	-- 0x25d3
		"11100111",	-- 0x25d4
		"01101101",	-- 0x25d5
		"11111011",	-- 0x25d6
		"00000001",	-- 0x25d7
		"01000100",	-- 0x25d8
		"00000001",	-- 0x25d9
		"11000101",	-- 0x25da
		"01001111",	-- 0x25db
		"01111100",	-- 0x25dc
		"10010010",	-- 0x25dd
		"01111011",	-- 0x25de
		"10110110",	-- 0x25df
		"00000001",	-- 0x25e0
		"00110011",	-- 0x25e1
		"10011010",	-- 0x25e2
		"01111000",	-- 0x25e3
		"01101110",	-- 0x25e4
		"10001111",	-- 0x25e5
		"00000000",	-- 0x25e6
		"01111000",	-- 0x25e7
		"11011011",	-- 0x25e8
		"01111010",	-- 0x25e9
		"00000001",	-- 0x25ea
		"11000101",	-- 0x25eb
		"01101101",	-- 0x25ec
		"01111110",	-- 0x25ed
		"01110000",	-- 0x25ee
		"01111011",	-- 0x25ef
		"01000110",	-- 0x25f0
		"11110010",	-- 0x25f1
		"01110101",	-- 0x25f2
		"00011000",	-- 0x25f3
		"10111000",	-- 0x25f4
		"00000001",	-- 0x25f5
		"00110101",	-- 0x25f6
		"01000100",	-- 0x25f7
		"00000011",	-- 0x25f8
		"00000001",	-- 0x25f9
		"11000100",	-- 0x25fa
		"11100111",	-- 0x25fb
		"01101000",	-- 0x25fc
		"11011010",	-- 0x25fd
		"01010000",	-- 0x25fe
		"11000100",	-- 0x25ff
		"01100001",	-- 0x2600
		"01000011",	-- 0x2601
		"00001110",	-- 0x2602
		"10001110",	-- 0x2603
		"00000000",	-- 0x2604
		"00000000",	-- 0x2605
		"00000001",	-- 0x2606
		"11000101",	-- 0x2607
		"01011011",	-- 0x2608
		"10000111",	-- 0x2609
		"00000001",	-- 0x260a
		"00000000",	-- 0x260b
		"01111110",	-- 0x260c
		"00000001",	-- 0x260d
		"11000101",	-- 0x260e
		"00000111",	-- 0x260f
		"01000001",	-- 0x2610
		"01111000",	-- 0x2611
		"00000001",	-- 0x2612
		"11000100",	-- 0x2613
		"11101001",	-- 0x2614
		"00110111",	-- 0x2615
		"00011000",	-- 0x2616
		"00001000",	-- 0x2617
		"10010111",	-- 0x2618
		"01010000",	-- 0x2619
		"01000101",	-- 0x261a
		"00001011",	-- 0x261b
		"01010010",	-- 0x261c
		"01010011",	-- 0x261d
		"01000000",	-- 0x261e
		"00000111",	-- 0x261f
		"10010111",	-- 0x2620
		"01010000",	-- 0x2621
		"01000100",	-- 0x2622
		"00000011",	-- 0x2623
		"10000110",	-- 0x2624
		"11111111",	-- 0x2625
		"11111111",	-- 0x2626
		"10111010",	-- 0x2627
		"00000010",	-- 0x2628
		"00001000",	-- 0x2629
		"10110110",	-- 0x262a
		"00000001",	-- 0x262b
		"00110001",	-- 0x262c
		"10111000",	-- 0x262d
		"00000001",	-- 0x262e
		"00110101",	-- 0x262f
		"01000101",	-- 0x2630
		"00000110",	-- 0x2631
		"01001010",	-- 0x2632
		"00001000",	-- 0x2633
		"11001010",	-- 0x2634
		"01111111",	-- 0x2635
		"01000000",	-- 0x2636
		"00000100",	-- 0x2637
		"01001011",	-- 0x2638
		"00000010",	-- 0x2639
		"11001010",	-- 0x263a
		"10000000",	-- 0x263b
		"10110010",	-- 0x263c
		"00000001",	-- 0x263d
		"01000110",	-- 0x263e
		"10110110",	-- 0x263f
		"00000001",	-- 0x2640
		"00110011",	-- 0x2641
		"10111000",	-- 0x2642
		"00000001",	-- 0x2643
		"00110101",	-- 0x2644
		"01000101",	-- 0x2645
		"00000110",	-- 0x2646
		"01001010",	-- 0x2647
		"00001000",	-- 0x2648
		"11001010",	-- 0x2649
		"01111111",	-- 0x264a
		"01000000",	-- 0x264b
		"00000100",	-- 0x264c
		"01001011",	-- 0x264d
		"00000010",	-- 0x264e
		"11001010",	-- 0x264f
		"10000000",	-- 0x2650
		"10110010",	-- 0x2651
		"00000001",	-- 0x2652
		"01000111",	-- 0x2653
		"00000001",	-- 0x2654
		"11101010",	-- 0x2655
		"00100010",	-- 0x2656
		"00000001",	-- 0x2657
		"11101000",	-- 0x2658
		"01100101",	-- 0x2659
		"11111010",	-- 0x265a
		"00000001",	-- 0x265b
		"11010110",	-- 0x265c
		"10010010",	-- 0x265d
		"01001110",	-- 0x265e
		"00110111",	-- 0x265f
		"00010110",	-- 0x2660
		"00000011",	-- 0x2661
		"00000011",	-- 0x2662
		"11100111",	-- 0x2663
		"01011110",	-- 0x2664
		"11001010",	-- 0x2665
		"01100001",	-- 0x2666
		"11010100",	-- 0x2667
		"10011000",	-- 0x2668
		"01000100",	-- 0x2669
		"00000001",	-- 0x266a
		"01010010",	-- 0x266b
		"10000001",	-- 0x266c
		"00010010",	-- 0x266d
		"01101000",	-- 0x266e
		"00000001",	-- 0x266f
		"11000100",	-- 0x2670
		"11011011",	-- 0x2671
		"10010011",	-- 0x2672
		"11111100",	-- 0x2673
		"01111000",	-- 0x2674
		"10110111",	-- 0x2675
		"00000010",	-- 0x2676
		"00001000",	-- 0x2677
		"01000100",	-- 0x2678
		"00000011",	-- 0x2679
		"10000110",	-- 0x267a
		"11111111",	-- 0x267b
		"11111111",	-- 0x267c
		"10001001",	-- 0x267d
		"00000000",	-- 0x267e
		"00000000",	-- 0x267f
		"01000100",	-- 0x2680
		"00000110",	-- 0x2681
		"10000110",	-- 0x2682
		"00000000",	-- 0x2683
		"00000000",	-- 0x2684
		"01110111",	-- 0x2685
		"01011000",	-- 0x2686
		"10001100",	-- 0x2687
		"01110101",	-- 0x2688
		"01011000",	-- 0x2689
		"00000001",	-- 0x268a
		"11000100",	-- 0x268b
		"11001100",	-- 0x268c
		"00111110",	-- 0x268d
		"01101110",	-- 0x268e
		"11111010",	-- 0x268f
		"00000001",	-- 0x2690
		"11001010",	-- 0x2691
		"00000001",	-- 0x2692
		"11000101",	-- 0x2693
		"01011011",	-- 0x2694
		"10001110",	-- 0x2695
		"01100100",	-- 0x2696
		"00000000",	-- 0x2697
		"00110101",	-- 0x2698
		"11010110",	-- 0x2699
		"00000011",	-- 0x269a
		"10001110",	-- 0x269b
		"01100100",	-- 0x269c
		"00000000",	-- 0x269d
		"00000001",	-- 0x269e
		"11000101",	-- 0x269f
		"10011011",	-- 0x26a0
		"10001000",	-- 0x26a1
		"00110011",	-- 0x26a2
		"00110011",	-- 0x26a3
		"01000100",	-- 0x26a4
		"00000010",	-- 0x26a5
		"01010010",	-- 0x26a6
		"01010011",	-- 0x26a7
		"10111010",	-- 0x26a8
		"00000001",	-- 0x26a9
		"11001000",	-- 0x26aa
		"01111110",	-- 0x26ab
		"10110110",	-- 0x26ac
		"00000001",	-- 0x26ad
		"00111000",	-- 0x26ae
		"00000001",	-- 0x26af
		"11000100",	-- 0x26b0
		"11001100",	-- 0x26b1
		"00000001",	-- 0x26b2
		"11000101",	-- 0x26b3
		"00000111",	-- 0x26b4
		"00110101",	-- 0x26b5
		"00010000",	-- 0x26b6
		"00010110",	-- 0x26b7
		"10011010",	-- 0x26b8
		"01111000",	-- 0x26b9
		"10110110",	-- 0x26ba
		"00000001",	-- 0x26bb
		"00100111",	-- 0x26bc
		"01001010",	-- 0x26bd
		"00001000",	-- 0x26be
		"10010111",	-- 0x26bf
		"01111000",	-- 0x26c0
		"01000101",	-- 0x26c1
		"00001011",	-- 0x26c2
		"01010010",	-- 0x26c3
		"01010011",	-- 0x26c4
		"01000000",	-- 0x26c5
		"00000111",	-- 0x26c6
		"10010111",	-- 0x26c7
		"01111000",	-- 0x26c8
		"01000100",	-- 0x26c9
		"00000011",	-- 0x26ca
		"10000110",	-- 0x26cb
		"11111111",	-- 0x26cc
		"11111111",	-- 0x26cd
		"10011010",	-- 0x26ce
		"01111000",	-- 0x26cf
		"01111001",	-- 0x26d0
		"00110000",	-- 0x26d1
		"01011001",	-- 0x26d2
		"01000100",	-- 0x26d3
		"00001000",	-- 0x26d4
		"01111001",	-- 0x26d5
		"00101100",	-- 0x26d6
		"01011001",	-- 0x26d7
		"01000100",	-- 0x26d8
		"00000101",	-- 0x26d9
		"01110101",	-- 0x26da
		"00111110",	-- 0x26db
		"10001100",	-- 0x26dc
		"01110111",	-- 0x26dd
		"00111110",	-- 0x26de
		"01111001",	-- 0x26df
		"00111001",	-- 0x26e0
		"01010000",	-- 0x26e1
		"01000101",	-- 0x26e2
		"00010000",	-- 0x26e3
		"00110101",	-- 0x26e4
		"01010110",	-- 0x26e5
		"00001101",	-- 0x26e6
		"01111001",	-- 0x26e7
		"11001010",	-- 0x26e8
		"01010111",	-- 0x26e9
		"01000101",	-- 0x26ea
		"00001000",	-- 0x26eb
		"01111001",	-- 0x26ec
		"11010010",	-- 0x26ed
		"01010111",	-- 0x26ee
		"01000101",	-- 0x26ef
		"00000101",	-- 0x26f0
		"01110111",	-- 0x26f1
		"00011110",	-- 0x26f2
		"10001100",	-- 0x26f3
		"01110101",	-- 0x26f4
		"00011110",	-- 0x26f5
		"10001111",	-- 0x26f6
		"00000001",	-- 0x26f7
		"00010010",	-- 0x26f8
		"10001110",	-- 0x26f9
		"11000010",	-- 0x26fa
		"01011011",	-- 0x26fb
		"00110111",	-- 0x26fc
		"00111110",	-- 0x26fd
		"00000011",	-- 0x26fe
		"10001110",	-- 0x26ff
		"11000010",	-- 0x2700
		"01011111",	-- 0x2701
		"01101110",	-- 0x2702
		"01101111",	-- 0x2703
		"11101010",	-- 0x2704
		"00000000",	-- 0x2705
		"10011110",	-- 0x2706
		"01111000",	-- 0x2707
		"00110101",	-- 0x2708
		"00010000",	-- 0x2709
		"00000011",	-- 0x270a
		"00110101",	-- 0x270b
		"00011110",	-- 0x270c
		"00000001",	-- 0x270d
		"01010010",	-- 0x270e
		"00000001",	-- 0x270f
		"11000101",	-- 0x2710
		"01011011",	-- 0x2711
		"10010111",	-- 0x2712
		"01111000",	-- 0x2713
		"01000100",	-- 0x2714
		"00000011",	-- 0x2715
		"10000110",	-- 0x2716
		"11111111",	-- 0x2717
		"11111111",	-- 0x2718
		"10001111",	-- 0x2719
		"11000011",	-- 0x271a
		"10111001",	-- 0x271b
		"00100001",	-- 0x271c
		"10100111",	-- 0x271d
		"01111111",	-- 0x271e
		"01111110",	-- 0x271f
		"10001010",	-- 0x2720
		"10001101",	-- 0x2721
		"00000001",	-- 0x2722
		"00011000",	-- 0x2723
		"01000010",	-- 0x2724
		"00000011",	-- 0x2725
		"00011100",	-- 0x2726
		"01000000",	-- 0x2727
		"11011001",	-- 0x2728
		"00110101",	-- 0x2729
		"11110110",	-- 0x272a
		"00000011",	-- 0x272b
		"00110111",	-- 0x272c
		"01111101",	-- 0x272d
		"00011011",	-- 0x272e
		"10000110",	-- 0x272f
		"00000010",	-- 0x2730
		"10010100",	-- 0x2731
		"00110101",	-- 0x2732
		"01010110",	-- 0x2733
		"00000011",	-- 0x2734
		"10000110",	-- 0x2735
		"00001010",	-- 0x2736
		"11001000",	-- 0x2737
		"00000101",	-- 0x2738
		"10111010",	-- 0x2739
		"00000001",	-- 0x273a
		"00001010",	-- 0x273b
		"10111010",	-- 0x273c
		"00000001",	-- 0x273d
		"00001100",	-- 0x273e
		"10111010",	-- 0x273f
		"00000001",	-- 0x2740
		"00001110",	-- 0x2741
		"10111010",	-- 0x2742
		"00000001",	-- 0x2743
		"00010000",	-- 0x2744
		"01110111",	-- 0x2745
		"11110101",	-- 0x2746
		"00000111",	-- 0x2747
		"01000000",	-- 0x2748
		"00010100",	-- 0x2749
		"10001110",	-- 0x274a
		"00000001",	-- 0x274b
		"00001010",	-- 0x274c
		"10001111",	-- 0x274d
		"00000001",	-- 0x274e
		"00010010",	-- 0x274f
		"00000101",	-- 0x2750
		"00011011",	-- 0x2751
		"10101010",	-- 0x2752
		"00000000",	-- 0x2753
		"00011100",	-- 0x2754
		"00011100",	-- 0x2755
		"10001100",	-- 0x2756
		"00000001",	-- 0x2757
		"00010000",	-- 0x2758
		"01000011",	-- 0x2759
		"11110110",	-- 0x275a
		"01110111",	-- 0x275b
		"11110101",	-- 0x275c
		"00000111",	-- 0x275d
		"11011010",	-- 0x275e
		"01001110",	-- 0x275f
		"10110010",	-- 0x2760
		"00000001",	-- 0x2761
		"11010110",	-- 0x2762
		"00000001",	-- 0x2763
		"11110011",	-- 0x2764
		"01110101",	-- 0x2765
		"01100011",	-- 0x2766
		"00000001",	-- 0x2767
		"11100101",	-- 0x2768
		"00111001",	-- 0x2769
		"00000100",	-- 0x276a
		"00000100",	-- 0x276b
		"00000100",	-- 0x276c
		"11001100",	-- 0x276d
		"00000101",	-- 0x276e
		"01000101",	-- 0x276f
		"00001010",	-- 0x2770
		"11000000",	-- 0x2771
		"00000101",	-- 0x2772
		"00000100",	-- 0x2773
		"11001100",	-- 0x2774
		"00001000",	-- 0x2775
		"01000101",	-- 0x2776
		"00000011",	-- 0x2777
		"11000000",	-- 0x2778
		"00001000",	-- 0x2779
		"00000100",	-- 0x277a
		"00111110",	-- 0x277b
		"10010110",	-- 0x277c
		"01011001",	-- 0x277d
		"00000100",	-- 0x277e
		"00000100",	-- 0x277f
		"11001100",	-- 0x2780
		"00000110",	-- 0x2781
		"01000101",	-- 0x2782
		"00000011",	-- 0x2783
		"11000000",	-- 0x2784
		"00000110",	-- 0x2785
		"00000100",	-- 0x2786
		"10001111",	-- 0x2787
		"11000000",	-- 0x2788
		"00000110",	-- 0x2789
		"00000001",	-- 0x278a
		"11000100",	-- 0x278b
		"10001010",	-- 0x278c
		"01101000",	-- 0x278d
		"00000001",	-- 0x278e
		"11000100",	-- 0x278f
		"11001101",	-- 0x2790
		"00111110",	-- 0x2791
		"10010110",	-- 0x2792
		"01011001",	-- 0x2793
		"10001111",	-- 0x2794
		"11000000",	-- 0x2795
		"11000111",	-- 0x2796
		"00000001",	-- 0x2797
		"11000100",	-- 0x2798
		"10000101",	-- 0x2799
		"10010010",	-- 0x279a
		"01111010",	-- 0x279b
		"01111110",	-- 0x279c
		"01100011",	-- 0x279d
		"10111110",	-- 0x279e
		"00000001",	-- 0x279f
		"00110001",	-- 0x27a0
		"00110111",	-- 0x27a1
		"00010110",	-- 0x27a2
		"00000011",	-- 0x27a3
		"00001010",	-- 0x27a4
		"00000001",	-- 0x27a5
		"00110011",	-- 0x27a6
		"10001111",	-- 0x27a7
		"00000001",	-- 0x27a8
		"00110011",	-- 0x27a9
		"11111011",	-- 0x27aa
		"00000001",	-- 0x27ab
		"00110111",	-- 0x27ac
		"00000001",	-- 0x27ad
		"11000101",	-- 0x27ae
		"01101101",	-- 0x27af
		"01100011",	-- 0x27b0
		"10110110",	-- 0x27b1
		"00000001",	-- 0x27b2
		"00110011",	-- 0x27b3
		"00110101",	-- 0x27b4
		"00010110",	-- 0x27b5
		"00010010",	-- 0x27b6
		"10111000",	-- 0x27b7
		"00000001",	-- 0x27b8
		"00110101",	-- 0x27b9
		"01000111",	-- 0x27ba
		"00010000",	-- 0x27bb
		"00010100",	-- 0x27bc
		"00010101",	-- 0x27bd
		"00011000",	-- 0x27be
		"00010101",	-- 0x27bf
		"10001001",	-- 0x27c0
		"00000000",	-- 0x27c1
		"00000000",	-- 0x27c2
		"01000110",	-- 0x27c3
		"00000001",	-- 0x27c4
		"01010111",	-- 0x27c5
		"10110111",	-- 0x27c6
		"00000001",	-- 0x27c7
		"00110101",	-- 0x27c8
		"10111010",	-- 0x27c9
		"00000001",	-- 0x27ca
		"00110101",	-- 0x27cb
		"01100011",	-- 0x27cc
		"10001111",	-- 0x27cd
		"11000001",	-- 0x27ce
		"01101000",	-- 0x27cf
		"11111011",	-- 0x27d0
		"00000001",	-- 0x27d1
		"00101001",	-- 0x27d2
		"01001010",	-- 0x27d3
		"00000011",	-- 0x27d4
		"10001111",	-- 0x27d5
		"11000001",	-- 0x27d6
		"01110010",	-- 0x27d7
		"10010110",	-- 0x27d8
		"01011001",	-- 0x27d9
		"00000001",	-- 0x27da
		"11000100",	-- 0x27db
		"00110000",	-- 0x27dc
		"10110010",	-- 0x27dd
		"00000001",	-- 0x27de
		"00111100",	-- 0x27df
		"00110101",	-- 0x27e0
		"10110100",	-- 0x27e1
		"00011010",	-- 0x27e2
		"10001111",	-- 0x27e3
		"11000001",	-- 0x27e4
		"10000101",	-- 0x27e5
		"00000001",	-- 0x27e6
		"11000100",	-- 0x27e7
		"01000010",	-- 0x27e8
		"01100001",	-- 0x27e9
		"01011000",	-- 0x27ea
		"10011010",	-- 0x27eb
		"01111000",	-- 0x27ec
		"10001111",	-- 0x27ed
		"11000001",	-- 0x27ee
		"01111100",	-- 0x27ef
		"00000001",	-- 0x27f0
		"11000100",	-- 0x27f1
		"01000010",	-- 0x27f2
		"10010111",	-- 0x27f3
		"01111000",	-- 0x27f4
		"01000100",	-- 0x27f5
		"00000011",	-- 0x27f6
		"10000110",	-- 0x27f7
		"11111111",	-- 0x27f8
		"11111111",	-- 0x27f9
		"10111010",	-- 0x27fa
		"00000001",	-- 0x27fb
		"00111101",	-- 0x27fc
		"10001111",	-- 0x27fd
		"11000001",	-- 0x27fe
		"10001110",	-- 0x27ff
		"00000001",	-- 0x2800
		"11000011",	-- 0x2801
		"11101110",	-- 0x2802
		"10011010",	-- 0x2803
		"01111000",	-- 0x2804
		"10001111",	-- 0x2805
		"11000001",	-- 0x2806
		"10110000",	-- 0x2807
		"00000001",	-- 0x2808
		"11000011",	-- 0x2809
		"11101110",	-- 0x280a
		"01100001",	-- 0x280b
		"00110110",	-- 0x280c
		"10110111",	-- 0x280d
		"00000001",	-- 0x280e
		"00111101",	-- 0x280f
		"01000100",	-- 0x2810
		"00000011",	-- 0x2811
		"10000110",	-- 0x2812
		"11111111",	-- 0x2813
		"11111111",	-- 0x2814
		"01100001",	-- 0x2815
		"00111000",	-- 0x2816
		"10111010",	-- 0x2817
		"00000001",	-- 0x2818
		"00111111",	-- 0x2819
		"10001111",	-- 0x281a
		"11000001",	-- 0x281b
		"10011111",	-- 0x281c
		"00000001",	-- 0x281d
		"11000011",	-- 0x281e
		"11101110",	-- 0x281f
		"10011010",	-- 0x2820
		"01111000",	-- 0x2821
		"10001111",	-- 0x2822
		"11000001",	-- 0x2823
		"11000001",	-- 0x2824
		"00000001",	-- 0x2825
		"11000011",	-- 0x2826
		"11101110",	-- 0x2827
		"01100001",	-- 0x2828
		"00011001",	-- 0x2829
		"01100001",	-- 0x282a
		"00100011",	-- 0x282b
		"10111010",	-- 0x282c
		"00000001",	-- 0x282d
		"01000001",	-- 0x282e
		"00000011",	-- 0x282f
		"11101010",	-- 0x2830
		"00010111",	-- 0x2831
		"00110111",	-- 0x2832
		"10110100",	-- 0x2833
		"00001101",	-- 0x2834
		"10110110",	-- 0x2835
		"00000001",	-- 0x2836
		"00111101",	-- 0x2837
		"10001000",	-- 0x2838
		"00000000",	-- 0x2839
		"00001100",	-- 0x283a
		"01000100",	-- 0x283b
		"00000010",	-- 0x283c
		"01010010",	-- 0x283d
		"01010011",	-- 0x283e
		"10111010",	-- 0x283f
		"00000001",	-- 0x2840
		"00111101",	-- 0x2841
		"01100011",	-- 0x2842
		"00111110",	-- 0x2843
		"11011010",	-- 0x2844
		"10010110",	-- 0x2845
		"00110101",	-- 0x2846
		"00010010",	-- 0x2847
		"00000010",	-- 0x2848
		"11001010",	-- 0x2849
		"00000000",	-- 0x284a
		"00000001",	-- 0x284b
		"11000101",	-- 0x284c
		"01011011",	-- 0x284d
		"01100011",	-- 0x284e
		"10010111",	-- 0x284f
		"01111000",	-- 0x2850
		"01000100",	-- 0x2851
		"00000011",	-- 0x2852
		"10000110",	-- 0x2853
		"11111111",	-- 0x2854
		"11111111",	-- 0x2855
		"00111110",	-- 0x2856
		"11111010",	-- 0x2857
		"00000010",	-- 0x2858
		"01000001",	-- 0x2859
		"00000001",	-- 0x285a
		"11000101",	-- 0x285b
		"01011011",	-- 0x285c
		"11000000",	-- 0x285d
		"00000100",	-- 0x285e
		"01000100",	-- 0x285f
		"00000011",	-- 0x2860
		"10000110",	-- 0x2861
		"11111111",	-- 0x2862
		"11111111",	-- 0x2863
		"01100011",	-- 0x2864
		"01110001",	-- 0x2865
		"01110001",	-- 0x2866
		"01000111",	-- 0x2867
		"00000011",	-- 0x2868
		"00000011",	-- 0x2869
		"11101010",	-- 0x286a
		"00001011",	-- 0x286b
		"10110110",	-- 0x286c
		"00000010",	-- 0x286d
		"00001000",	-- 0x286e
		"10001111",	-- 0x286f
		"11000001",	-- 0x2870
		"01010100",	-- 0x2871
		"00000001",	-- 0x2872
		"11000100",	-- 0x2873
		"00110000",	-- 0x2874
		"00000100",	-- 0x2875
		"00110101",	-- 0x2876
		"10110100",	-- 0x2877
		"00010111",	-- 0x2878
		"10111010",	-- 0x2879
		"00000001",	-- 0x287a
		"00101011",	-- 0x287b
		"10111010",	-- 0x287c
		"00000001",	-- 0x287d
		"00101101",	-- 0x287e
		"10111010",	-- 0x287f
		"00000001",	-- 0x2880
		"00101111",	-- 0x2881
		"01010010",	-- 0x2882
		"01010011",	-- 0x2883
		"10111010",	-- 0x2884
		"00000001",	-- 0x2885
		"00101001",	-- 0x2886
		"10111010",	-- 0x2887
		"00000001",	-- 0x2888
		"00100111",	-- 0x2889
		"00110011",	-- 0x288a
		"11111111",	-- 0x288b
		"10101010",	-- 0x288c
		"00000011",	-- 0x288d
		"11101010",	-- 0x288e
		"00001011",	-- 0x288f
		"01101000",	-- 0x2890
		"10111110",	-- 0x2891
		"00000001",	-- 0x2892
		"00101111",	-- 0x2893
		"10111001",	-- 0x2894
		"00000001",	-- 0x2895
		"00101111",	-- 0x2896
		"01000100",	-- 0x2897
		"00000100",	-- 0x2898
		"00111110",	-- 0x2899
		"10110110",	-- 0x289a
		"00000001",	-- 0x289b
		"00101111",	-- 0x289c
		"10011010",	-- 0x289d
		"01111000",	-- 0x289e
		"00111010",	-- 0x289f
		"01111010",	-- 0x28a0
		"10001111",	-- 0x28a1
		"00000000",	-- 0x28a2
		"01111000",	-- 0x28a3
		"10110110",	-- 0x28a4
		"00000001",	-- 0x28a5
		"00101011",	-- 0x28a6
		"00000001",	-- 0x28a7
		"11000011",	-- 0x28a8
		"11100000",	-- 0x28a9
		"01101000",	-- 0x28aa
		"01110101",	-- 0x28ab
		"00011000",	-- 0x28ac
		"10111000",	-- 0x28ad
		"00000001",	-- 0x28ae
		"00101011",	-- 0x28af
		"01000100",	-- 0x28b0
		"00000011",	-- 0x28b1
		"00000001",	-- 0x28b2
		"11000100",	-- 0x28b3
		"11100111",	-- 0x28b4
		"10001001",	-- 0x28b5
		"00000001",	-- 0x28b6
		"00000000",	-- 0x28b7
		"01000101",	-- 0x28b8
		"00101001",	-- 0x28b9
		"00111110",	-- 0x28ba
		"11111010",	-- 0x28bb
		"00000010",	-- 0x28bc
		"01000000",	-- 0x28bd
		"00110111",	-- 0x28be
		"00011000",	-- 0x28bf
		"00000011",	-- 0x28c0
		"11111010",	-- 0x28c1
		"00000010",	-- 0x28c2
		"00111111",	-- 0x28c3
		"01010100",	-- 0x28c4
		"11001100",	-- 0x28c5
		"00000000",	-- 0x28c6
		"01000110",	-- 0x28c7
		"00000001",	-- 0x28c8
		"01010000",	-- 0x28c9
		"10000001",	-- 0x28ca
		"10000000",	-- 0x28cb
		"00000001",	-- 0x28cc
		"11000101",	-- 0x28cd
		"00000111",	-- 0x28ce
		"00111100",	-- 0x28cf
		"00000001",	-- 0x28d0
		"11000100",	-- 0x28d1
		"11101001",	-- 0x28d2
		"10110111",	-- 0x28d3
		"00000001",	-- 0x28d4
		"00101001",	-- 0x28d5
		"01001000",	-- 0x28d6
		"00001000",	-- 0x28d7
		"10000110",	-- 0x28d8
		"01111111",	-- 0x28d9
		"11111111",	-- 0x28da
		"00110111",	-- 0x28db
		"00011000",	-- 0x28dc
		"00000010",	-- 0x28dd
		"01010110",	-- 0x28de
		"01010111",	-- 0x28df
		"10111010",	-- 0x28e0
		"00000001",	-- 0x28e1
		"00101001",	-- 0x28e2
		"01111000",	-- 0x28e3
		"10111010",	-- 0x28e4
		"00000001",	-- 0x28e5
		"00101011",	-- 0x28e6
		"10001111",	-- 0x28e7
		"00000000",	-- 0x28e8
		"01111000",	-- 0x28e9
		"10110110",	-- 0x28ea
		"00000001",	-- 0x28eb
		"00101101",	-- 0x28ec
		"00000001",	-- 0x28ed
		"11000011",	-- 0x28ee
		"11100000",	-- 0x28ef
		"10111010",	-- 0x28f0
		"00000001",	-- 0x28f1
		"00101101",	-- 0x28f2
		"01111000",	-- 0x28f3
		"00111111",	-- 0x28f4
		"00110111",	-- 0x28f5
		"00010011",	-- 0x28f6
		"00000010",	-- 0x28f7
		"01110010",	-- 0x28f8
		"10101010",	-- 0x28f9
		"01111001",	-- 0x28fa
		"00000010",	-- 0x28fb
		"10101010",	-- 0x28fc
		"01000100",	-- 0x28fd
		"00001000",	-- 0x28fe
		"01110110",	-- 0x28ff
		"10101010",	-- 0x2900
		"00110101",	-- 0x2901
		"01010110",	-- 0x2902
		"00000011",	-- 0x2903
		"10000111",	-- 0x2904
		"00000001",	-- 0x2905
		"11110100",	-- 0x2906
		"10111000",	-- 0x2907
		"00000001",	-- 0x2908
		"00101101",	-- 0x2909
		"10111110",	-- 0x290a
		"00000001",	-- 0x290b
		"00101101",	-- 0x290c
		"00001010",	-- 0x290d
		"00000001",	-- 0x290e
		"00101111",	-- 0x290f
		"10111110",	-- 0x2910
		"00000001",	-- 0x2911
		"00101011",	-- 0x2912
		"00001010",	-- 0x2913
		"00000001",	-- 0x2914
		"00101101",	-- 0x2915
		"01101001",	-- 0x2916
		"00001010",	-- 0x2917
		"00000001",	-- 0x2918
		"00101011",	-- 0x2919
		"01110101",	-- 0x291a
		"00011000",	-- 0x291b
		"01000100",	-- 0x291c
		"00000011",	-- 0x291d
		"00000001",	-- 0x291e
		"11000100",	-- 0x291f
		"11100111",	-- 0x2920
		"00111110",	-- 0x2921
		"11111011",	-- 0x2922
		"00000010",	-- 0x2923
		"00111101",	-- 0x2924
		"00110111",	-- 0x2925
		"00011000",	-- 0x2926
		"00000011",	-- 0x2927
		"11111011",	-- 0x2928
		"00000010",	-- 0x2929
		"00111110",	-- 0x292a
		"00000001",	-- 0x292b
		"11000101",	-- 0x292c
		"01001111",	-- 0x292d
		"10011010",	-- 0x292e
		"01111000",	-- 0x292f
		"10001111",	-- 0x2930
		"11000001",	-- 0x2931
		"01100011",	-- 0x2932
		"00000001",	-- 0x2933
		"11000100",	-- 0x2934
		"00110111",	-- 0x2935
		"10010010",	-- 0x2936
		"01111010",	-- 0x2937
		"11111010",	-- 0x2938
		"00000010",	-- 0x2939
		"00111111",	-- 0x293a
		"00110111",	-- 0x293b
		"00011000",	-- 0x293c
		"00000011",	-- 0x293d
		"11111010",	-- 0x293e
		"00000010",	-- 0x293f
		"01000000",	-- 0x2940
		"10010001",	-- 0x2941
		"01111010",	-- 0x2942
		"00000110",	-- 0x2943
		"01000100",	-- 0x2944
		"00000010",	-- 0x2945
		"11001010",	-- 0x2946
		"11111111",	-- 0x2947
		"01011011",	-- 0x2948
		"01010101",	-- 0x2949
		"11001101",	-- 0x294a
		"00000000",	-- 0x294b
		"01000110",	-- 0x294c
		"00000001",	-- 0x294d
		"01010001",	-- 0x294e
		"01101101",	-- 0x294f
		"10011110",	-- 0x2950
		"01111000",	-- 0x2951
		"00000001",	-- 0x2952
		"11000101",	-- 0x2953
		"01011011",	-- 0x2954
		"01011000",	-- 0x2955
		"01001010",	-- 0x2956
		"00000011",	-- 0x2957
		"10000110",	-- 0x2958
		"01111111",	-- 0x2959
		"11111111",	-- 0x295a
		"00000001",	-- 0x295b
		"11000100",	-- 0x295c
		"11101001",	-- 0x295d
		"10011010",	-- 0x295e
		"01111010",	-- 0x295f
		"10011110",	-- 0x2960
		"01111000",	-- 0x2961
		"01111100",	-- 0x2962
		"10000001",	-- 0x2963
		"10000000",	-- 0x2964
		"00000001",	-- 0x2965
		"11000101",	-- 0x2966
		"00000111",	-- 0x2967
		"00111100",	-- 0x2968
		"00000001",	-- 0x2969
		"11000100",	-- 0x296a
		"11101001",	-- 0x296b
		"10011010",	-- 0x296c
		"01111000",	-- 0x296d
		"01110101",	-- 0x296e
		"00011000",	-- 0x296f
		"10110110",	-- 0x2970
		"00000001",	-- 0x2971
		"00101001",	-- 0x2972
		"01001010",	-- 0x2973
		"00000011",	-- 0x2974
		"00000001",	-- 0x2975
		"11000100",	-- 0x2976
		"11100111",	-- 0x2977
		"00111110",	-- 0x2978
		"01101000",	-- 0x2979
		"11111010",	-- 0x297a
		"00000001",	-- 0x297b
		"00111100",	-- 0x297c
		"01101100",	-- 0x297d
		"10000001",	-- 0x297e
		"10000000",	-- 0x297f
		"00000100",	-- 0x2980
		"00000100",	-- 0x2981
		"01010100",	-- 0x2982
		"01010101",	-- 0x2983
		"10000100",	-- 0x2984
		"00000000",	-- 0x2985
		"10001001",	-- 0x2986
		"00000000",	-- 0x2987
		"00000000",	-- 0x2988
		"01000110",	-- 0x2989
		"00000010",	-- 0x298a
		"01010000",	-- 0x298b
		"01010001",	-- 0x298c
		"00000001",	-- 0x298d
		"11000101",	-- 0x298e
		"00000111",	-- 0x298f
		"00111100",	-- 0x2990
		"00000001",	-- 0x2991
		"11000100",	-- 0x2992
		"11101001",	-- 0x2993
		"10010111",	-- 0x2994
		"01111000",	-- 0x2995
		"01001000",	-- 0x2996
		"00001000",	-- 0x2997
		"10000110",	-- 0x2998
		"01111111",	-- 0x2999
		"11111111",	-- 0x299a
		"00110111",	-- 0x299b
		"00011000",	-- 0x299c
		"00000010",	-- 0x299d
		"01010110",	-- 0x299e
		"01010111",	-- 0x299f
		"00000001",	-- 0x29a0
		"11101010",	-- 0x29a1
		"00001100",	-- 0x29a2
		"10111010",	-- 0x29a3
		"00000001",	-- 0x29a4
		"00101001",	-- 0x29a5
		"01111100",	-- 0x29a6
		"01111110",	-- 0x29a7
		"00000001",	-- 0x29a8
		"11000101",	-- 0x29a9
		"01011011",	-- 0x29aa
		"00000100",	-- 0x29ab
		"00000100",	-- 0x29ac
		"00000001",	-- 0x29ad
		"11000100",	-- 0x29ae
		"11101001",	-- 0x29af
		"10010111",	-- 0x29b0
		"01111010",	-- 0x29b1
		"01001000",	-- 0x29b2
		"00001000",	-- 0x29b3
		"10000110",	-- 0x29b4
		"01111111",	-- 0x29b5
		"11111111",	-- 0x29b6
		"00110111",	-- 0x29b7
		"00011000",	-- 0x29b8
		"00000010",	-- 0x29b9
		"01010110",	-- 0x29ba
		"01010111",	-- 0x29bb
		"00000001",	-- 0x29bc
		"11101010",	-- 0x29bd
		"00001100",	-- 0x29be
		"00111110",	-- 0x29bf
		"01110101",	-- 0x29c0
		"00011000",	-- 0x29c1
		"01011000",	-- 0x29c2
		"01001010",	-- 0x29c3
		"00000011",	-- 0x29c4
		"00000001",	-- 0x29c5
		"11000100",	-- 0x29c6
		"11100111",	-- 0x29c7
		"01101000",	-- 0x29c8
		"10001001",	-- 0x29c9
		"00000000",	-- 0x29ca
		"00100000",	-- 0x29cb
		"01000100",	-- 0x29cc
		"00100010",	-- 0x29cd
		"10000110",	-- 0x29ce
		"00000000",	-- 0x29cf
		"01000000",	-- 0x29d0
		"10010010",	-- 0x29d1
		"01111001",	-- 0x29d2
		"10010011",	-- 0x29d3
		"01111011",	-- 0x29d4
		"11111010",	-- 0x29d5
		"00000001",	-- 0x29d6
		"01000001",	-- 0x29d7
		"10010010",	-- 0x29d8
		"01111010",	-- 0x29d9
		"11111010",	-- 0x29da
		"00000001",	-- 0x29db
		"00111111",	-- 0x29dc
		"10010010",	-- 0x29dd
		"01111100",	-- 0x29de
		"00110011",	-- 0x29df
		"00000010",	-- 0x29e0
		"01111000",	-- 0x29e1
		"00111100",	-- 0x29e2
		"10000111",	-- 0x29e3
		"00000000",	-- 0x29e4
		"00100000",	-- 0x29e5
		"01011010",	-- 0x29e6
		"01010011",	-- 0x29e7
		"10001111",	-- 0x29e8
		"00000000",	-- 0x29e9
		"01111000",	-- 0x29ea
		"00000001",	-- 0x29eb
		"11000011",	-- 0x29ec
		"11110100",	-- 0x29ed
		"01000000",	-- 0x29ee
		"00001001",	-- 0x29ef
		"10110110",	-- 0x29f0
		"00000001",	-- 0x29f1
		"00111111",	-- 0x29f2
		"00110111",	-- 0x29f3
		"00011000",	-- 0x29f4
		"00000011",	-- 0x29f5
		"10110110",	-- 0x29f6
		"00000001",	-- 0x29f7
		"01000001",	-- 0x29f8
		"00111110",	-- 0x29f9
		"01111000",	-- 0x29fa
		"00000110",	-- 0x29fb
		"00000001",	-- 0x29fc
		"11000101",	-- 0x29fd
		"00000111",	-- 0x29fe
		"00000001",	-- 0x29ff
		"11000101",	-- 0x2a00
		"00111001",	-- 0x2a01
		"00000001",	-- 0x2a02
		"11000100",	-- 0x2a03
		"11101001",	-- 0x2a04
		"10111010",	-- 0x2a05
		"00000001",	-- 0x2a06
		"00100111",	-- 0x2a07
		"00000001",	-- 0x2a08
		"11101000",	-- 0x2a09
		"00110010",	-- 0x2a0a
		"01100011",	-- 0x2a0b
		"01011000",	-- 0x2a0c
		"01001010",	-- 0x2a0d
		"00000111",	-- 0x2a0e
		"01111001",	-- 0x2a0f
		"01111010",	-- 0x2a10
		"11010000",	-- 0x2a11
		"01000100",	-- 0x2a12
		"00000010",	-- 0x2a13
		"01010010",	-- 0x2a14
		"01010011",	-- 0x2a15
		"01100011",	-- 0x2a16
		"01100001",	-- 0x2a17
		"00001001",	-- 0x2a18
		"00000001",	-- 0x2a19
		"11101000",	-- 0x2a1a
		"01100101",	-- 0x2a1b
		"00000000",	-- 0x2a1c
		"00000000",	-- 0x2a1d
		"00000000",	-- 0x2a1e
		"00000011",	-- 0x2a1f
		"11000111",	-- 0x2a20
		"01001001",	-- 0x2a21
		"01111001",	-- 0x2a22
		"00111101",	-- 0x2a23
		"11000111",	-- 0x2a24
		"01000101",	-- 0x2a25
		"00000110",	-- 0x2a26
		"01110111",	-- 0x2a27
		"01010101",	-- 0x2a28
		"01110101",	-- 0x2a29
		"10010101",	-- 0x2a2a
		"01110101",	-- 0x2a2b
		"00010101",	-- 0x2a2c
		"10001111",	-- 0x2a2d
		"11000010",	-- 0x2a2e
		"01100111",	-- 0x2a2f
		"11011010",	-- 0x2a30
		"01010110",	-- 0x2a31
		"01010011",	-- 0x2a32
		"00000001",	-- 0x2a33
		"11000011",	-- 0x2a34
		"11110100",	-- 0x2a35
		"10010010",	-- 0x2a36
		"01111000",	-- 0x2a37
		"10001111",	-- 0x2a38
		"11000010",	-- 0x2a39
		"01110010",	-- 0x2a3a
		"00000001",	-- 0x2a3b
		"11000011",	-- 0x2a3c
		"11110010",	-- 0x2a3d
		"10010001",	-- 0x2a3e
		"01111000",	-- 0x2a3f
		"00000001",	-- 0x2a40
		"11000100",	-- 0x2a41
		"11001011",	-- 0x2a42
		"10111010",	-- 0x2a43
		"00000001",	-- 0x2a44
		"01110011",	-- 0x2a45
		"10001111",	-- 0x2a46
		"11000010",	-- 0x2a47
		"01111101",	-- 0x2a48
		"00000001",	-- 0x2a49
		"11000011",	-- 0x2a4a
		"11110010",	-- 0x2a4b
		"10110010",	-- 0x2a4c
		"00000001",	-- 0x2a4d
		"01110010",	-- 0x2a4e
		"11111010",	-- 0x2a4f
		"00000001",	-- 0x2a50
		"11010010",	-- 0x2a51
		"10010010",	-- 0x2a52
		"01001110",	-- 0x2a53
		"10001111",	-- 0x2a54
		"11000010",	-- 0x2a55
		"11110010",	-- 0x2a56
		"11011011",	-- 0x2a57
		"01011011",	-- 0x2a58
		"00000001",	-- 0x2a59
		"11000100",	-- 0x2a5a
		"01000100",	-- 0x2a5b
		"10010010",	-- 0x2a5c
		"01111010",	-- 0x2a5d
		"00110101",	-- 0x2a5e
		"01010110",	-- 0x2a5f
		"00001001",	-- 0x2a60
		"11111010",	-- 0x2a61
		"00000001",	-- 0x2a62
		"00110011",	-- 0x2a63
		"11000000",	-- 0x2a64
		"00001010",	-- 0x2a65
		"11011100",	-- 0x2a66
		"01111010",	-- 0x2a67
		"01000100",	-- 0x2a68
		"00000100",	-- 0x2a69
		"01110111",	-- 0x2a6a
		"00011110",	-- 0x2a6b
		"01110010",	-- 0x2a6c
		"10100011",	-- 0x2a6d
		"01111001",	-- 0x2a6e
		"11010010",	-- 0x2a6f
		"01010111",	-- 0x2a70
		"01000101",	-- 0x2a71
		"00000101",	-- 0x2a72
		"01111001",	-- 0x2a73
		"01111000",	-- 0x2a74
		"01011011",	-- 0x2a75
		"01000101",	-- 0x2a76
		"00000010",	-- 0x2a77
		"01110101",	-- 0x2a78
		"00011110",	-- 0x2a79
		"00110111",	-- 0x2a7a
		"00011110",	-- 0x2a7b
		"00011000",	-- 0x2a7c
		"11111011",	-- 0x2a7d
		"00000001",	-- 0x2a7e
		"01000111",	-- 0x2a7f
		"11001101",	-- 0x2a80
		"00000110",	-- 0x2a81
		"01001101",	-- 0x2a82
		"00010001",	-- 0x2a83
		"11111010",	-- 0x2a84
		"00000001",	-- 0x2a85
		"00110011",	-- 0x2a86
		"11011100",	-- 0x2a87
		"01111010",	-- 0x2a88
		"01000101",	-- 0x2a89
		"00001010",	-- 0x2a8a
		"10001111",	-- 0x2a8b
		"11000010",	-- 0x2a8c
		"11110111",	-- 0x2a8d
		"00000001",	-- 0x2a8e
		"11000011",	-- 0x2a8f
		"11110010",	-- 0x2a90
		"10010010",	-- 0x2a91
		"10100011",	-- 0x2a92
		"01110101",	-- 0x2a93
		"00011110",	-- 0x2a94
		"01000000",	-- 0x2a95
		"00010101",	-- 0x2a96
		"11011010",	-- 0x2a97
		"10100011",	-- 0x2a98
		"01000111",	-- 0x2a99
		"00000111",	-- 0x2a9a
		"11000100",	-- 0x2a9b
		"00001001",	-- 0x2a9c
		"01000100",	-- 0x2a9d
		"00000001",	-- 0x2a9e
		"01010010",	-- 0x2a9f
		"10010010",	-- 0x2aa0
		"10100011",	-- 0x2aa1
		"01100011",	-- 0x2aa2
		"11011010",	-- 0x2aa3
		"10100011",	-- 0x2aa4
		"11001100",	-- 0x2aa5
		"00101011",	-- 0x2aa6
		"01000011",	-- 0x2aa7
		"00000010",	-- 0x2aa8
		"11001010",	-- 0x2aa9
		"00101011",	-- 0x2aaa
		"01100011",	-- 0x2aab
		"11011010",	-- 0x2aac
		"01001110",	-- 0x2aad
		"10110010",	-- 0x2aae
		"00000001",	-- 0x2aaf
		"11010010",	-- 0x2ab0
		"11111010",	-- 0x2ab1
		"00000001",	-- 0x2ab2
		"11010011",	-- 0x2ab3
		"10010010",	-- 0x2ab4
		"01001110",	-- 0x2ab5
		"00110101",	-- 0x2ab6
		"11010000",	-- 0x2ab7
		"00100111",	-- 0x2ab8
		"01111001",	-- 0x2ab9
		"01011100",	-- 0x2aba
		"11010000",	-- 0x2abb
		"01000101",	-- 0x2abc
		"00100010",	-- 0x2abd
		"11011011",	-- 0x2abe
		"11111011",	-- 0x2abf
		"10001111",	-- 0x2ac0
		"11000010",	-- 0x2ac1
		"11001101",	-- 0x2ac2
		"00000001",	-- 0x2ac3
		"11000100",	-- 0x2ac4
		"01000100",	-- 0x2ac5
		"11011100",	-- 0x2ac6
		"01011011",	-- 0x2ac7
		"01000011",	-- 0x2ac8
		"00010110",	-- 0x2ac9
		"01111001",	-- 0x2aca
		"00101000",	-- 0x2acb
		"01011011",	-- 0x2acc
		"01000101",	-- 0x2acd
		"00010001",	-- 0x2ace
		"01111001",	-- 0x2acf
		"00000011",	-- 0x2ad0
		"01011101",	-- 0x2ad1
		"01000101",	-- 0x2ad2
		"00001100",	-- 0x2ad3
		"01111001",	-- 0x2ad4
		"11010010",	-- 0x2ad5
		"01010111",	-- 0x2ad6
		"01000101",	-- 0x2ad7
		"00000111",	-- 0x2ad8
		"01111001",	-- 0x2ad9
		"10010011",	-- 0x2ada
		"01010110",	-- 0x2adb
		"01000101",	-- 0x2adc
		"00000010",	-- 0x2add
		"01110111",	-- 0x2ade
		"00111110",	-- 0x2adf
		"11111010",	-- 0x2ae0
		"00000001",	-- 0x2ae1
		"01000111",	-- 0x2ae2
		"11111011",	-- 0x2ae3
		"00000001",	-- 0x2ae4
		"00110011",	-- 0x2ae5
		"10011010",	-- 0x2ae6
		"01111000",	-- 0x2ae7
		"00110111",	-- 0x2ae8
		"01010110",	-- 0x2ae9
		"00000100",	-- 0x2aea
		"01110010",	-- 0x2aeb
		"11011001",	-- 0x2aec
		"01110101",	-- 0x2aed
		"00111110",	-- 0x2aee
		"00110111",	-- 0x2aef
		"00111001",	-- 0x2af0
		"00000110",	-- 0x2af1
		"01110101",	-- 0x2af2
		"00011110",	-- 0x2af3
		"01110101",	-- 0x2af4
		"01011110",	-- 0x2af5
		"01000000",	-- 0x2af6
		"00111010",	-- 0x2af7
		"11001100",	-- 0x2af8
		"11111110",	-- 0x2af9
		"01001101",	-- 0x2afa
		"00111011",	-- 0x2afb
		"00110101",	-- 0x2afc
		"01011110",	-- 0x2afd
		"00001100",	-- 0x2afe
		"11001100",	-- 0x2aff
		"00000101",	-- 0x2b00
		"01001101",	-- 0x2b01
		"00001000",	-- 0x2b02
		"11001101",	-- 0x2b03
		"00100001",	-- 0x2b04
		"01000101",	-- 0x2b05
		"00000100",	-- 0x2b06
		"01110010",	-- 0x2b07
		"10111101",	-- 0x2b08
		"01110111",	-- 0x2b09
		"01011110",	-- 0x2b0a
		"10001111",	-- 0x2b0b
		"11000010",	-- 0x2b0c
		"11100111",	-- 0x2b0d
		"11011011",	-- 0x2b0e
		"11111011",	-- 0x2b0f
		"00000001",	-- 0x2b10
		"11000100",	-- 0x2b11
		"01000100",	-- 0x2b12
		"11011100",	-- 0x2b13
		"10111101",	-- 0x2b14
		"01000101",	-- 0x2b15
		"00100000",	-- 0x2b16
		"10010110",	-- 0x2b17
		"01111000",	-- 0x2b18
		"00110111",	-- 0x2b19
		"00111110",	-- 0x2b1a
		"00011101",	-- 0x2b1b
		"00110101",	-- 0x2b1c
		"00011110",	-- 0x2b1d
		"00011010",	-- 0x2b1e
		"11001100",	-- 0x2b1f
		"00001001",	-- 0x2b20
		"01001101",	-- 0x2b21
		"00010110",	-- 0x2b22
		"11001101",	-- 0x2b23
		"01001101",	-- 0x2b24
		"01000101",	-- 0x2b25
		"00010010",	-- 0x2b26
		"01111001",	-- 0x2b27
		"00011111",	-- 0x2b28
		"11011001",	-- 0x2b29
		"01000100",	-- 0x2b2a
		"00001101",	-- 0x2b2b
		"01110111",	-- 0x2b2c
		"01111110",	-- 0x2b2d
		"01110111",	-- 0x2b2e
		"00011110",	-- 0x2b2f
		"01000000",	-- 0x2b30
		"00000111",	-- 0x2b31
		"11001010",	-- 0x2b32
		"11111111",	-- 0x2b33
		"10110010",	-- 0x2b34
		"00000001",	-- 0x2b35
		"01011110",	-- 0x2b36
		"01110101",	-- 0x2b37
		"01111110",	-- 0x2b38
		"10010110",	-- 0x2b39
		"01111000",	-- 0x2b3a
		"00110111",	-- 0x2b3b
		"00010100",	-- 0x2b3c
		"00000011",	-- 0x2b3d
		"00110111",	-- 0x2b3e
		"01010110",	-- 0x2b3f
		"00001000",	-- 0x2b40
		"11001100",	-- 0x2b41
		"00001000",	-- 0x2b42
		"01001101",	-- 0x2b43
		"00001111",	-- 0x2b44
		"11001101",	-- 0x2b45
		"00100110",	-- 0x2b46
		"01000101",	-- 0x2b47
		"00001011",	-- 0x2b48
		"01010010",	-- 0x2b49
		"10010010",	-- 0x2b4a
		"11011010",	-- 0x2b4b
		"10110010",	-- 0x2b4c
		"00000001",	-- 0x2b4d
		"01100010",	-- 0x2b4e
		"11011010",	-- 0x2b4f
		"01011011",	-- 0x2b50
		"10110010",	-- 0x2b51
		"00000001",	-- 0x2b52
		"01100111",	-- 0x2b53
		"00000011",	-- 0x2b54
		"11101100",	-- 0x2b55
		"00100100",	-- 0x2b56
		"00110111",	-- 0x2b57
		"01111110",	-- 0x2b58
		"00001100",	-- 0x2b59
		"11111011",	-- 0x2b5a
		"00000001",	-- 0x2b5b
		"01010111",	-- 0x2b5c
		"10001111",	-- 0x2b5d
		"11000010",	-- 0x2b5e
		"11010100",	-- 0x2b5f
		"00000001",	-- 0x2b60
		"11000100",	-- 0x2b61
		"01000100",	-- 0x2b62
		"10110010",	-- 0x2b63
		"00000001",	-- 0x2b64
		"01011110",	-- 0x2b65
		"10010110",	-- 0x2b66
		"01011001",	-- 0x2b67
		"10001001",	-- 0x2b68
		"01010100",	-- 0x2b69
		"00000000",	-- 0x2b6a
		"01000100",	-- 0x2b6b
		"00000011",	-- 0x2b6c
		"00000001",	-- 0x2b6d
		"11001000",	-- 0x2b6e
		"11000000",	-- 0x2b6f
		"10111010",	-- 0x2b70
		"00000001",	-- 0x2b71
		"01100011",	-- 0x2b72
		"00111110",	-- 0x2b73
		"10111000",	-- 0x2b74
		"00000001",	-- 0x2b75
		"01100101",	-- 0x2b76
		"01000101",	-- 0x2b77
		"00000101",	-- 0x2b78
		"00000001",	-- 0x2b79
		"11000100",	-- 0x2b7a
		"11100000",	-- 0x2b7b
		"01000000",	-- 0x2b7c
		"00000110",	-- 0x2b7d
		"01010011",	-- 0x2b7e
		"11011010",	-- 0x2b7f
		"01011011",	-- 0x2b80
		"10110010",	-- 0x2b81
		"00000001",	-- 0x2b82
		"01100111",	-- 0x2b83
		"10110011",	-- 0x2b84
		"00000001",	-- 0x2b85
		"01100001",	-- 0x2b86
		"00001010",	-- 0x2b87
		"00000001",	-- 0x2b88
		"01100101",	-- 0x2b89
		"00110101",	-- 0x2b8a
		"01010110",	-- 0x2b8b
		"00011110",	-- 0x2b8c
		"11011010",	-- 0x2b8d
		"01011011",	-- 0x2b8e
		"11110100",	-- 0x2b8f
		"00000001",	-- 0x2b90
		"01100111",	-- 0x2b91
		"01000100",	-- 0x2b92
		"00000001",	-- 0x2b93
		"01010010",	-- 0x2b94
		"11001100",	-- 0x2b95
		"00001110",	-- 0x2b96
		"01000100",	-- 0x2b97
		"00010010",	-- 0x2b98
		"00110111",	-- 0x2b99
		"00111110",	-- 0x2b9a
		"00001111",	-- 0x2b9b
		"11011010",	-- 0x2b9c
		"11111011",	-- 0x2b9d
		"11001100",	-- 0x2b9e
		"00100000",	-- 0x2b9f
		"01000101",	-- 0x2ba0
		"00001001",	-- 0x2ba1
		"11001100",	-- 0x2ba2
		"10001101",	-- 0x2ba3
		"01000100",	-- 0x2ba4
		"00000101",	-- 0x2ba5
		"01111001",	-- 0x2ba6
		"10011001",	-- 0x2ba7
		"11011001",	-- 0x2ba8
		"01000101",	-- 0x2ba9
		"00001000",	-- 0x2baa
		"10000110",	-- 0x2bab
		"11111111",	-- 0x2bac
		"11111110",	-- 0x2bad
		"10110010",	-- 0x2bae
		"00000001",	-- 0x2baf
		"01100010",	-- 0x2bb0
		"10010011",	-- 0x2bb1
		"11011010",	-- 0x2bb2
		"11111011",	-- 0x2bb3
		"00000001",	-- 0x2bb4
		"01100001",	-- 0x2bb5
		"11110101",	-- 0x2bb6
		"00000001",	-- 0x2bb7
		"01100010",	-- 0x2bb8
		"01000100",	-- 0x2bb9
		"00000001",	-- 0x2bba
		"01010011",	-- 0x2bbb
		"10001111",	-- 0x2bbc
		"11000010",	-- 0x2bbd
		"11011011",	-- 0x2bbe
		"00000001",	-- 0x2bbf
		"11000100",	-- 0x2bc0
		"01000100",	-- 0x2bc1
		"01101000",	-- 0x2bc2
		"10001111",	-- 0x2bc3
		"11000010",	-- 0x2bc4
		"11101110",	-- 0x2bc5
		"11011011",	-- 0x2bc6
		"01010010",	-- 0x2bc7
		"00000001",	-- 0x2bc8
		"11000100",	-- 0x2bc9
		"00111110",	-- 0x2bca
		"01011011",	-- 0x2bcb
		"01111110",	-- 0x2bcc
		"00000001",	-- 0x2bcd
		"11000101",	-- 0x2bce
		"01001111",	-- 0x2bcf
		"11110100",	-- 0x2bd0
		"00000001",	-- 0x2bd1
		"01010111",	-- 0x2bd2
		"01000101",	-- 0x2bd3
		"00000001",	-- 0x2bd4
		"01010010",	-- 0x2bd5
		"01010100",	-- 0x2bd6
		"10110010",	-- 0x2bd7
		"00000001",	-- 0x2bd8
		"01011111",	-- 0x2bd9
		"11111100",	-- 0x2bda
		"00000001",	-- 0x2bdb
		"01011110",	-- 0x2bdc
		"01000011",	-- 0x2bdd
		"00000011",	-- 0x2bde
		"11111010",	-- 0x2bdf
		"00000001",	-- 0x2be0
		"01011110",	-- 0x2be1
		"11110000",	-- 0x2be2
		"00000001",	-- 0x2be3
		"01100000",	-- 0x2be4
		"01000100",	-- 0x2be5
		"00000010",	-- 0x2be6
		"11001010",	-- 0x2be7
		"11111111",	-- 0x2be8
		"11001100",	-- 0x2be9
		"00000000",	-- 0x2bea
		"01000100",	-- 0x2beb
		"00000010",	-- 0x2bec
		"11001010",	-- 0x2bed
		"00000000",	-- 0x2bee
		"10110010",	-- 0x2bef
		"00000001",	-- 0x2bf0
		"01011101",	-- 0x2bf1
		"01100011",	-- 0x2bf2
		"11111011",	-- 0x2bf3
		"00000001",	-- 0x2bf4
		"11010011",	-- 0x2bf5
		"11001111",	-- 0x2bf6
		"00001000",	-- 0x2bf7
		"01000110",	-- 0x2bf8
		"00001100",	-- 0x2bf9
		"11001011",	-- 0x2bfa
		"00000100",	-- 0x2bfb
		"11110001",	-- 0x2bfc
		"00000001",	-- 0x2bfd
		"01011110",	-- 0x2bfe
		"01000100",	-- 0x2bff
		"00000010",	-- 0x2c00
		"11001011",	-- 0x2c01
		"11111111",	-- 0x2c02
		"10110011",	-- 0x2c03
		"00000001",	-- 0x2c04
		"01011110",	-- 0x2c05
		"01100011",	-- 0x2c06
		"01010010",	-- 0x2c07
		"01111001",	-- 0x2c08
		"00010100",	-- 0x2c09
		"11011010",	-- 0x2c0a
		"01000101",	-- 0x2c0b
		"00001001",	-- 0x2c0c
		"11111010",	-- 0x2c0d
		"00000001",	-- 0x2c0e
		"01100010",	-- 0x2c0f
		"11000000",	-- 0x2c10
		"00000100",	-- 0x2c11
		"01000100",	-- 0x2c12
		"00000010",	-- 0x2c13
		"11001010",	-- 0x2c14
		"11111111",	-- 0x2c15
		"10110010",	-- 0x2c16
		"00000001",	-- 0x2c17
		"01100010",	-- 0x2c18
		"01100011",	-- 0x2c19
		"10001111",	-- 0x2c1a
		"11000010",	-- 0x2c1b
		"11100010",	-- 0x2c1c
		"00000001",	-- 0x2c1d
		"11000011",	-- 0x2c1e
		"11101110",	-- 0x2c1f
		"10110010",	-- 0x2c20
		"00000001",	-- 0x2c21
		"01100000",	-- 0x2c22
		"01100011",	-- 0x2c23
		"11011010",	-- 0x2c24
		"01001110",	-- 0x2c25
		"10110010",	-- 0x2c26
		"00000001",	-- 0x2c27
		"11010011",	-- 0x2c28
		"00000001",	-- 0x2c29
		"11110110",	-- 0x2c2a
		"11000101",	-- 0x2c2b
		"01110001",	-- 0x2c2c
		"00110001",	-- 0x2c2d
		"01000111",	-- 0x2c2e
		"00000011",	-- 0x2c2f
		"00000011",	-- 0x2c30
		"11101111",	-- 0x2c31
		"10110000",	-- 0x2c32
		"00000001",	-- 0x2c33
		"11101010",	-- 0x2c34
		"10010111",	-- 0x2c35
		"11011010",	-- 0x2c36
		"01010111",	-- 0x2c37
		"01111001",	-- 0x2c38
		"00110010",	-- 0x2c39
		"01011001",	-- 0x2c3a
		"01000101",	-- 0x2c3b
		"00000100",	-- 0x2c3c
		"11001100",	-- 0x2c3d
		"10000110",	-- 0x2c3e
		"01000100",	-- 0x2c3f
		"00001100",	-- 0x2c40
		"11001100",	-- 0x2c41
		"11011100",	-- 0x2c42
		"01000100",	-- 0x2c43
		"00001000",	-- 0x2c44
		"00110101",	-- 0x2c45
		"01010110",	-- 0x2c46
		"01000010",	-- 0x2c47
		"01111001",	-- 0x2c48
		"01100001",	-- 0x2c49
		"01010000",	-- 0x2c4a
		"01000011",	-- 0x2c4b
		"00010101",	-- 0x2c4c
		"11111010",	-- 0x2c4d
		"00000001",	-- 0x2c4e
		"01010110",	-- 0x2c4f
		"11000100",	-- 0x2c50
		"10000000",	-- 0x2c51
		"01000111",	-- 0x2c52
		"00111101",	-- 0x2c53
		"01000010",	-- 0x2c54
		"00000100",	-- 0x2c55
		"11000000",	-- 0x2c56
		"00000001",	-- 0x2c57
		"01000000",	-- 0x2c58
		"00000010",	-- 0x2c59
		"11000100",	-- 0x2c5a
		"00000001",	-- 0x2c5b
		"01000101",	-- 0x2c5c
		"00110011",	-- 0x2c5d
		"11000000",	-- 0x2c5e
		"10000000",	-- 0x2c5f
		"01000000",	-- 0x2c60
		"00110001",	-- 0x2c61
		"10010010",	-- 0x2c62
		"01111000",	-- 0x2c63
		"10001111",	-- 0x2c64
		"11000010",	-- 0x2c65
		"10000100",	-- 0x2c66
		"00000001",	-- 0x2c67
		"11000011",	-- 0x2c68
		"11110000",	-- 0x2c69
		"10010010",	-- 0x2c6a
		"01111100",	-- 0x2c6b
		"11011010",	-- 0x2c6c
		"01111000",	-- 0x2c6d
		"10001111",	-- 0x2c6e
		"11000010",	-- 0x2c6f
		"10010101",	-- 0x2c70
		"00000001",	-- 0x2c71
		"11000011",	-- 0x2c72
		"11110000",	-- 0x2c73
		"10010010",	-- 0x2c74
		"01111010",	-- 0x2c75
		"10000110",	-- 0x2c76
		"01001110",	-- 0x2c77
		"01010111",	-- 0x2c78
		"10010010",	-- 0x2c79
		"01111001",	-- 0x2c7a
		"10010011",	-- 0x2c7b
		"01111011",	-- 0x2c7c
		"00110011",	-- 0x2c7d
		"00000010",	-- 0x2c7e
		"01111000",	-- 0x2c7f
		"10010110",	-- 0x2c80
		"01010000",	-- 0x2c81
		"10001111",	-- 0x2c82
		"00000000",	-- 0x2c83
		"01111000",	-- 0x2c84
		"00000001",	-- 0x2c85
		"11000011",	-- 0x2c86
		"11110100",	-- 0x2c87
		"01000000",	-- 0x2c88
		"00001001",	-- 0x2c89
		"10001111",	-- 0x2c8a
		"11000010",	-- 0x2c8b
		"10100110",	-- 0x2c8c
		"00000001",	-- 0x2c8d
		"11000011",	-- 0x2c8e
		"11110000",	-- 0x2c8f
		"10001100",	-- 0x2c90
		"11001010",	-- 0x2c91
		"10000000",	-- 0x2c92
		"10110010",	-- 0x2c93
		"00000001",	-- 0x2c94
		"01010110",	-- 0x2c95
		"11111010",	-- 0x2c96
		"00000001",	-- 0x2c97
		"11010100",	-- 0x2c98
		"10010010",	-- 0x2c99
		"01001110",	-- 0x2c9a
		"11001010",	-- 0x2c9b
		"01010101",	-- 0x2c9c
		"00110111",	-- 0x2c9d
		"01010110",	-- 0x2c9e
		"00011110",	-- 0x2c9f
		"01111001",	-- 0x2ca0
		"01011100",	-- 0x2ca1
		"11010000",	-- 0x2ca2
		"01000101",	-- 0x2ca3
		"00011001",	-- 0x2ca4
		"01111001",	-- 0x2ca5
		"00111101",	-- 0x2ca6
		"11010010",	-- 0x2ca7
		"01000101",	-- 0x2ca8
		"00010100",	-- 0x2ca9
		"10010110",	-- 0x2caa
		"01110100",	-- 0x2cab
		"10000111",	-- 0x2cac
		"00000000",	-- 0x2cad
		"11000000",	-- 0x2cae
		"10011000",	-- 0x2caf
		"01011001",	-- 0x2cb0
		"01000100",	-- 0x2cb1
		"00000010",	-- 0x2cb2
		"01010010",	-- 0x2cb3
		"01010011",	-- 0x2cb4
		"00000001",	-- 0x2cb5
		"11000100",	-- 0x2cb6
		"11100000",	-- 0x2cb7
		"10001111",	-- 0x2cb8
		"11000010",	-- 0x2cb9
		"10110111",	-- 0x2cba
		"00000001",	-- 0x2cbb
		"11000100",	-- 0x2cbc
		"01000100",	-- 0x2cbd
		"10010010",	-- 0x2cbe
		"01111000",	-- 0x2cbf
		"01110101",	-- 0x2cc0
		"00011110",	-- 0x2cc1
		"00110101",	-- 0x2cc2
		"11010110",	-- 0x2cc3
		"00000111",	-- 0x2cc4
		"00110111",	-- 0x2cc5
		"00111110",	-- 0x2cc6
		"00001010",	-- 0x2cc7
		"01110101",	-- 0x2cc8
		"00111110",	-- 0x2cc9
		"01000000",	-- 0x2cca
		"00000100",	-- 0x2ccb
		"01110001",	-- 0x2ccc
		"00111110",	-- 0x2ccd
		"01000110",	-- 0x2cce
		"00000010",	-- 0x2ccf
		"01110111",	-- 0x2cd0
		"00011110",	-- 0x2cd1
		"00110101",	-- 0x2cd2
		"11010010",	-- 0x2cd3
		"00000111",	-- 0x2cd4
		"00110111",	-- 0x2cd5
		"01011110",	-- 0x2cd6
		"00001010",	-- 0x2cd7
		"01110101",	-- 0x2cd8
		"01011110",	-- 0x2cd9
		"01000000",	-- 0x2cda
		"00000100",	-- 0x2cdb
		"01110001",	-- 0x2cdc
		"01011110",	-- 0x2cdd
		"01000110",	-- 0x2cde
		"00000010",	-- 0x2cdf
		"01110111",	-- 0x2ce0
		"00011110",	-- 0x2ce1
		"00110101",	-- 0x2ce2
		"00010110",	-- 0x2ce3
		"00011100",	-- 0x2ce4
		"00110111",	-- 0x2ce5
		"01010110",	-- 0x2ce6
		"00100001",	-- 0x2ce7
		"01111001",	-- 0x2ce8
		"00101000",	-- 0x2ce9
		"01011011",	-- 0x2cea
		"01000100",	-- 0x2ceb
		"00011100",	-- 0x2cec
		"01111001",	-- 0x2ced
		"00010101",	-- 0x2cee
		"01011011",	-- 0x2cef
		"01000101",	-- 0x2cf0
		"00010111",	-- 0x2cf1
		"01111001",	-- 0x2cf2
		"00000010",	-- 0x2cf3
		"01011101",	-- 0x2cf4
		"01000100",	-- 0x2cf5
		"00010010",	-- 0x2cf6
		"01111001",	-- 0x2cf7
		"11100100",	-- 0x2cf8
		"01010111",	-- 0x2cf9
		"01000101",	-- 0x2cfa
		"00001101",	-- 0x2cfb
		"00110101",	-- 0x2cfc
		"00011110",	-- 0x2cfd
		"00001010",	-- 0x2cfe
		"01000000",	-- 0x2cff
		"00100010",	-- 0x2d00
		"01010010",	-- 0x2d01
		"01010011",	-- 0x2d02
		"10111010",	-- 0x2d03
		"00000001",	-- 0x2d04
		"01111111",	-- 0x2d05
		"10111010",	-- 0x2d06
		"00000001",	-- 0x2d07
		"10000001",	-- 0x2d08
		"01110010",	-- 0x2d09
		"11011000",	-- 0x2d0a
		"01100001",	-- 0x2d0b
		"00001100",	-- 0x2d0c
		"01100001",	-- 0x2d0d
		"00000011",	-- 0x2d0e
		"00000011",	-- 0x2d0f
		"11101101",	-- 0x2d10
		"01101110",	-- 0x2d11
		"00000101",	-- 0x2d12
		"01010010",	-- 0x2d13
		"10110010",	-- 0x2d14
		"00000001",	-- 0x2d15
		"01111000",	-- 0x2d16
		"00000111",	-- 0x2d17
		"01100011",	-- 0x2d18
		"10000110",	-- 0x2d19
		"10000000",	-- 0x2d1a
		"10000000",	-- 0x2d1b
		"10111010",	-- 0x2d1c
		"00000001",	-- 0x2d1d
		"01111011",	-- 0x2d1e
		"10111010",	-- 0x2d1f
		"00000001",	-- 0x2d20
		"01111101",	-- 0x2d21
		"01100011",	-- 0x2d22
		"11111010",	-- 0x2d23
		"00000001",	-- 0x2d24
		"01111000",	-- 0x2d25
		"11001100",	-- 0x2d26
		"00100000",	-- 0x2d27
		"01000101",	-- 0x2d28
		"01000100",	-- 0x2d29
		"01100001",	-- 0x2d2a
		"11100110",	-- 0x2d2b
		"10001111",	-- 0x2d2c
		"00000001",	-- 0x2d2d
		"01111011",	-- 0x2d2e
		"01101111",	-- 0x2d2f
		"01111110",	-- 0x2d30
		"00011101",	-- 0x2d31
		"10001101",	-- 0x2d32
		"00000001",	-- 0x2d33
		"01111111",	-- 0x2d34
		"01000100",	-- 0x2d35
		"00001000",	-- 0x2d36
		"11101010",	-- 0x2d37
		"00000000",	-- 0x2d38
		"11101100",	-- 0x2d39
		"10000000",	-- 0x2d3a
		"01000100",	-- 0x2d3b
		"11110100",	-- 0x2d3c
		"01000000",	-- 0x2d3d
		"11110000",	-- 0x2d3e
		"11101010",	-- 0x2d3f
		"00000000",	-- 0x2d40
		"11001100",	-- 0x2d41
		"10000011",	-- 0x2d42
		"01000101",	-- 0x2d43
		"00001110",	-- 0x2d44
		"11101010",	-- 0x2d45
		"00000100",	-- 0x2d46
		"11000000",	-- 0x2d47
		"00001001",	-- 0x2d48
		"11001100",	-- 0x2d49
		"00110011",	-- 0x2d4a
		"01000011",	-- 0x2d4b
		"00000010",	-- 0x2d4c
		"11001010",	-- 0x2d4d
		"00110011",	-- 0x2d4e
		"10100010",	-- 0x2d4f
		"00000100",	-- 0x2d50
		"01100001",	-- 0x2d51
		"11000110",	-- 0x2d52
		"10001111",	-- 0x2d53
		"00000001",	-- 0x2d54
		"01111111",	-- 0x2d55
		"00011010",	-- 0x2d56
		"01000111",	-- 0x2d57
		"00010101",	-- 0x2d58
		"10001101",	-- 0x2d59
		"00000001",	-- 0x2d5a
		"10000011",	-- 0x2d5b
		"01000101",	-- 0x2d5c
		"11111000",	-- 0x2d5d
		"10001111",	-- 0x2d5e
		"00000001",	-- 0x2d5f
		"01111111",	-- 0x2d60
		"11101010",	-- 0x2d61
		"10000000",	-- 0x2d62
		"11000100",	-- 0x2d63
		"00001001",	-- 0x2d64
		"01000100",	-- 0x2d65
		"00000001",	-- 0x2d66
		"01010010",	-- 0x2d67
		"10000010",	-- 0x2d68
		"10001101",	-- 0x2d69
		"00000001",	-- 0x2d6a
		"10000011",	-- 0x2d6b
		"01000101",	-- 0x2d6c
		"11110011",	-- 0x2d6d
		"11011010",	-- 0x2d6e
		"11011000",	-- 0x2d6f
		"01000110",	-- 0x2d70
		"00010011",	-- 0x2d71
		"00000101",	-- 0x2d72
		"10001111",	-- 0x2d73
		"00000001",	-- 0x2d74
		"01111111",	-- 0x2d75
		"11001010",	-- 0x2d76
		"00101011",	-- 0x2d77
		"11101100",	-- 0x2d78
		"10000000",	-- 0x2d79
		"01000100",	-- 0x2d7a
		"00000010",	-- 0x2d7b
		"10100010",	-- 0x2d7c
		"10000000",	-- 0x2d7d
		"00011101",	-- 0x2d7e
		"10001101",	-- 0x2d7f
		"00000001",	-- 0x2d80
		"10000011",	-- 0x2d81
		"01000101",	-- 0x2d82
		"11110100",	-- 0x2d83
		"00000111",	-- 0x2d84
		"11011011",	-- 0x2d85
		"01111000",	-- 0x2d86
		"01111001",	-- 0x2d87
		"00000110",	-- 0x2d88
		"11011000",	-- 0x2d89
		"01000101",	-- 0x2d8a
		"00110101",	-- 0x2d8b
		"01010010",	-- 0x2d8c
		"01010011",	-- 0x2d8d
		"10001111",	-- 0x2d8e
		"00000001",	-- 0x2d8f
		"01111111",	-- 0x2d90
		"11100001",	-- 0x2d91
		"10000000",	-- 0x2d92
		"10000000",	-- 0x2d93
		"00000000",	-- 0x2d94
		"00011101",	-- 0x2d95
		"10001101",	-- 0x2d96
		"00000001",	-- 0x2d97
		"10000011",	-- 0x2d98
		"01000101",	-- 0x2d99
		"11110110",	-- 0x2d9a
		"00000001",	-- 0x2d9b
		"11000100",	-- 0x2d9c
		"11011111",	-- 0x2d9d
		"10010011",	-- 0x2d9e
		"01111001",	-- 0x2d9f
		"11011011",	-- 0x2da0
		"10100001",	-- 0x2da1
		"00010001",	-- 0x2da2
		"00010001",	-- 0x2da3
		"00010001",	-- 0x2da4
		"00010001",	-- 0x2da5
		"11000001",	-- 0x2da6
		"00000010",	-- 0x2da7
		"11000011",	-- 0x2da8
		"00000011",	-- 0x2da9
		"10001111",	-- 0x2daa
		"00000001",	-- 0x2dab
		"01111111",	-- 0x2dac
		"00001111",	-- 0x2dad
		"01010010",	-- 0x2dae
		"11011011",	-- 0x2daf
		"01111000",	-- 0x2db0
		"11100001",	-- 0x2db1
		"10000000",	-- 0x2db2
		"10000000",	-- 0x2db3
		"00000000",	-- 0x2db4
		"11010101",	-- 0x2db5
		"01111001",	-- 0x2db6
		"10000100",	-- 0x2db7
		"00000000",	-- 0x2db8
		"01000111",	-- 0x2db9
		"00000110",	-- 0x2dba
		"01000101",	-- 0x2dbb
		"00000011",	-- 0x2dbc
		"11001011",	-- 0x2dbd
		"11111111",	-- 0x2dbe
		"01000001",	-- 0x2dbf
		"01010011",	-- 0x2dc0
		"10001111",	-- 0x2dc1
		"11000011",	-- 0x2dc2
		"10111111",	-- 0x2dc3
		"00100001",	-- 0x2dc4
		"10011000",	-- 0x2dc5
		"10110011",	-- 0x2dc6
		"00000001",	-- 0x2dc7
		"01011000",	-- 0x2dc8
		"01000000",	-- 0x2dc9
		"01010010",	-- 0x2dca
		"01111001",	-- 0x2dcb
		"01011100",	-- 0x2dcc
		"11011000",	-- 0x2dcd
		"01000101",	-- 0x2dce
		"00110011",	-- 0x2dcf
		"10001110",	-- 0x2dd0
		"00000001",	-- 0x2dd1
		"01111011",	-- 0x2dd2
		"11011010",	-- 0x2dd3
		"10100010",	-- 0x2dd4
		"00010000",	-- 0x2dd5
		"00010000",	-- 0x2dd6
		"00010000",	-- 0x2dd7
		"00010000",	-- 0x2dd8
		"11000010",	-- 0x2dd9
		"00000011",	-- 0x2dda
		"00001100",	-- 0x2ddb
		"11101010",	-- 0x2ddc
		"00000000",	-- 0x2ddd
		"10000001",	-- 0x2dde
		"00000111",	-- 0x2ddf
		"01101000",	-- 0x2de0
		"10010110",	-- 0x2de1
		"11110110",	-- 0x2de2
		"10111000",	-- 0x2de3
		"00000001",	-- 0x2de4
		"01111001",	-- 0x2de5
		"01111111",	-- 0x2de6
		"10000111",	-- 0x2de7
		"00000100",	-- 0x2de8
		"00100100",	-- 0x2de9
		"01001010",	-- 0x2dea
		"00000010",	-- 0x2deb
		"01010010",	-- 0x2dec
		"01010011",	-- 0x2ded
		"00000001",	-- 0x2dee
		"11000100",	-- 0x2def
		"11011110",	-- 0x2df0
		"11001101",	-- 0x2df1
		"10110011",	-- 0x2df2
		"01000101",	-- 0x2df3
		"00010100",	-- 0x2df4
		"11101010",	-- 0x2df5
		"00000100",	-- 0x2df6
		"01000111",	-- 0x2df7
		"00000111",	-- 0x2df8
		"11000100",	-- 0x2df9
		"00011010",	-- 0x2dfa
		"01000100",	-- 0x2dfb
		"00000001",	-- 0x2dfc
		"01010010",	-- 0x2dfd
		"10100010",	-- 0x2dfe
		"00000100",	-- 0x2dff
		"00000001",	-- 0x2e00
		"11101101",	-- 0x2e01
		"00011001",	-- 0x2e02
		"01010010",	-- 0x2e03
		"10110010",	-- 0x2e04
		"00000001",	-- 0x2e05
		"01111000",	-- 0x2e06
		"01000000",	-- 0x2e07
		"00000111",	-- 0x2e08
		"00001111",	-- 0x2e09
		"00111101",	-- 0x2e0a
		"00000001",	-- 0x2e0b
		"11000100",	-- 0x2e0c
		"11011110",	-- 0x2e0d
		"10100011",	-- 0x2e0e
		"00000000",	-- 0x2e0f
		"10010110",	-- 0x2e10
		"11110110",	-- 0x2e11
		"10111010",	-- 0x2e12
		"00000001",	-- 0x2e13
		"01111001",	-- 0x2e14
		"11111010",	-- 0x2e15
		"00000001",	-- 0x2e16
		"01111000",	-- 0x2e17
		"01010110",	-- 0x2e18
		"10110010",	-- 0x2e19
		"00000001",	-- 0x2e1a
		"01111000",	-- 0x2e1b
		"01100011",	-- 0x2e1c
		"11011010",	-- 0x2e1d
		"01001110",	-- 0x2e1e
		"10110010",	-- 0x2e1f
		"00000001",	-- 0x2e20
		"11010100",	-- 0x2e21
		"11111010",	-- 0x2e22
		"00000010",	-- 0x2e23
		"00111100",	-- 0x2e24
		"00110111",	-- 0x2e25
		"01010110",	-- 0x2e26
		"00110111",	-- 0x2e27
		"01011011",	-- 0x2e28
		"01010010",	-- 0x2e29
		"00000110",	-- 0x2e2a
		"10000111",	-- 0x2e2b
		"00000000",	-- 0x2e2c
		"01010101",	-- 0x2e2d
		"11110101",	-- 0x2e2e
		"00000001",	-- 0x2e2f
		"01011000",	-- 0x2e30
		"10000100",	-- 0x2e31
		"00000000",	-- 0x2e32
		"01000100",	-- 0x2e33
		"00000010",	-- 0x2e34
		"01010010",	-- 0x2e35
		"01010011",	-- 0x2e36
		"00000001",	-- 0x2e37
		"11000100",	-- 0x2e38
		"11100000",	-- 0x2e39
		"10010011",	-- 0x2e3a
		"01111000",	-- 0x2e3b
		"10001111",	-- 0x2e3c
		"11000010",	-- 0x2e3d
		"11000000",	-- 0x2e3e
		"11011011",	-- 0x2e3f
		"01011011",	-- 0x2e40
		"00000001",	-- 0x2e41
		"11000100",	-- 0x2e42
		"01000111",	-- 0x2e43
		"10001110",	-- 0x2e44
		"11000010",	-- 0x2e45
		"11001001",	-- 0x2e46
		"00110111",	-- 0x2e47
		"11010110",	-- 0x2e48
		"00000001",	-- 0x2e49
		"00011100",	-- 0x2e4a
		"00110101",	-- 0x2e4b
		"11010010",	-- 0x2e4c
		"00000010",	-- 0x2e4d
		"00011100",	-- 0x2e4e
		"00011100",	-- 0x2e4f
		"11101100",	-- 0x2e50
		"00000000",	-- 0x2e51
		"01000100",	-- 0x2e52
		"00000010",	-- 0x2e53
		"11101010",	-- 0x2e54
		"00000000",	-- 0x2e55
		"11011100",	-- 0x2e56
		"01111000",	-- 0x2e57
		"01000011",	-- 0x2e58
		"00000101",	-- 0x2e59
		"00000001",	-- 0x2e5a
		"11101101",	-- 0x2e5b
		"00010010",	-- 0x2e5c
		"11011010",	-- 0x2e5d
		"01111000",	-- 0x2e5e
		"10110010",	-- 0x2e5f
		"00000001",	-- 0x2e60
		"01010101",	-- 0x2e61
		"11111011",	-- 0x2e62
		"00000001",	-- 0x2e63
		"01011100",	-- 0x2e64
		"11011010",	-- 0x2e65
		"10100110",	-- 0x2e66
		"11001100",	-- 0x2e67
		"11111111",	-- 0x2e68
		"01000111",	-- 0x2e69
		"00011011",	-- 0x2e6a
		"01011000",	-- 0x2e6b
		"01000110",	-- 0x2e6c
		"00001010",	-- 0x2e6d
		"11001011",	-- 0x2e6e
		"00101011",	-- 0x2e6f
		"00110101",	-- 0x2e70
		"01010011",	-- 0x2e71
		"00011011",	-- 0x2e72
		"00110101",	-- 0x2e73
		"01110011",	-- 0x2e74
		"00011000",	-- 0x2e75
		"01000000",	-- 0x2e76
		"00010001",	-- 0x2e77
		"11001100",	-- 0x2e78
		"00001100",	-- 0x2e79
		"01000100",	-- 0x2e7a
		"00000110",	-- 0x2e7b
		"11000101",	-- 0x2e7c
		"00000001",	-- 0x2e7d
		"01000100",	-- 0x2e7e
		"00001001",	-- 0x2e7f
		"01000000",	-- 0x2e80
		"00000100",	-- 0x2e81
		"11000101",	-- 0x2e82
		"00001001",	-- 0x2e83
		"01000100",	-- 0x2e84
		"00000011",	-- 0x2e85
		"01010011",	-- 0x2e86
		"11001010",	-- 0x2e87
		"11111110",	-- 0x2e88
		"01010110",	-- 0x2e89
		"01000111",	-- 0x2e8a
		"00000010",	-- 0x2e8b
		"10010010",	-- 0x2e8c
		"10100110",	-- 0x2e8d
		"10110011",	-- 0x2e8e
		"00000001",	-- 0x2e8f
		"01011100",	-- 0x2e90
		"01000000",	-- 0x2e91
		"00101010",	-- 0x2e92
		"00110111",	-- 0x2e93
		"01110011",	-- 0x2e94
		"00010001",	-- 0x2e95
		"01111001",	-- 0x2e96
		"00001010",	-- 0x2e97
		"01011101",	-- 0x2e98
		"01000101",	-- 0x2e99
		"00001001",	-- 0x2e9a
		"01111001",	-- 0x2e9b
		"00101001",	-- 0x2e9c
		"01010010",	-- 0x2e9d
		"01000101",	-- 0x2e9e
		"00000100",	-- 0x2e9f
		"01110010",	-- 0x2ea0
		"10100110",	-- 0x2ea1
		"01000000",	-- 0x2ea2
		"00000011",	-- 0x2ea3
		"00110011",	-- 0x2ea4
		"11111111",	-- 0x2ea5
		"10100110",	-- 0x2ea6
		"01100011",	-- 0x2ea7
		"00110111",	-- 0x2ea8
		"01010011",	-- 0x2ea9
		"00010001",	-- 0x2eaa
		"01111001",	-- 0x2eab
		"00001010",	-- 0x2eac
		"01011101",	-- 0x2ead
		"01000101",	-- 0x2eae
		"00001001",	-- 0x2eaf
		"01111001",	-- 0x2eb0
		"00101001",	-- 0x2eb1
		"01010010",	-- 0x2eb2
		"01000101",	-- 0x2eb3
		"00000100",	-- 0x2eb4
		"01110010",	-- 0x2eb5
		"10100110",	-- 0x2eb6
		"01000000",	-- 0x2eb7
		"00000011",	-- 0x2eb8
		"00110011",	-- 0x2eb9
		"11111111",	-- 0x2eba
		"10100110",	-- 0x2ebb
		"01100011",	-- 0x2ebc
		"00000001",	-- 0x2ebd
		"11101010",	-- 0x2ebe
		"10100011",	-- 0x2ebf
		"11110000",	-- 0x2ec0
		"00000010",	-- 0x2ec1
		"00010110",	-- 0x2ec2
		"01000100",	-- 0x2ec3
		"00000010",	-- 0x2ec4
		"11001010",	-- 0x2ec5
		"11111111",	-- 0x2ec6
		"11111011",	-- 0x2ec7
		"00000010",	-- 0x2ec8
		"01000011",	-- 0x2ec9
		"11001111",	-- 0x2eca
		"00001111",	-- 0x2ecb
		"01000111",	-- 0x2ecc
		"00000110",	-- 0x2ecd
		"11000000",	-- 0x2ece
		"00011010",	-- 0x2ecf
		"01000100",	-- 0x2ed0
		"00000010",	-- 0x2ed1
		"11001010",	-- 0x2ed2
		"11111111",	-- 0x2ed3
		"11110000",	-- 0x2ed4
		"00000001",	-- 0x2ed5
		"01011100",	-- 0x2ed6
		"01000100",	-- 0x2ed7
		"00000010",	-- 0x2ed8
		"11001010",	-- 0x2ed9
		"11111111",	-- 0x2eda
		"10110010",	-- 0x2edb
		"00000010",	-- 0x2edc
		"00011011",	-- 0x2edd
		"11111010",	-- 0x2ede
		"00000001",	-- 0x2edf
		"11010101",	-- 0x2ee0
		"10010010",	-- 0x2ee1
		"01001110",	-- 0x2ee2
		"01111001",	-- 0x2ee3
		"10000111",	-- 0x2ee4
		"01011100",	-- 0x2ee5
		"01000010",	-- 0x2ee6
		"00000101",	-- 0x2ee7
		"01111001",	-- 0x2ee8
		"00100100",	-- 0x2ee9
		"01011011",	-- 0x2eea
		"01000100",	-- 0x2eeb
		"00000100",	-- 0x2eec
		"01110101",	-- 0x2eed
		"11011110",	-- 0x2eee
		"01000000",	-- 0x2eef
		"00110100",	-- 0x2ef0
		"00110101",	-- 0x2ef1
		"11010000",	-- 0x2ef2
		"00110001",	-- 0x2ef3
		"00110111",	-- 0x2ef4
		"11011110",	-- 0x2ef5
		"00000111",	-- 0x2ef6
		"01110101",	-- 0x2ef7
		"11011110",	-- 0x2ef8
		"10000110",	-- 0x2ef9
		"00000000",	-- 0x2efa
		"00000000",	-- 0x2efb
		"01000000",	-- 0x2efc
		"00101001",	-- 0x2efd
		"10110110",	-- 0x2efe
		"00000001",	-- 0x2eff
		"01011010",	-- 0x2f00
		"11001100",	-- 0x2f01
		"11111110",	-- 0x2f02
		"01000100",	-- 0x2f03
		"00100000",	-- 0x2f04
		"00110101",	-- 0x2f05
		"01010110",	-- 0x2f06
		"00001111",	-- 0x2f07
		"10001001",	-- 0x2f08
		"00000000",	-- 0x2f09
		"01010110",	-- 0x2f0a
		"01000101",	-- 0x2f0b
		"00000101",	-- 0x2f0c
		"10000111",	-- 0x2f0d
		"00000000",	-- 0x2f0e
		"00001001",	-- 0x2f0f
		"01000000",	-- 0x2f10
		"00010101",	-- 0x2f11
		"10000111",	-- 0x2f12
		"00000000",	-- 0x2f13
		"00100010",	-- 0x2f14
		"01000000",	-- 0x2f15
		"00010000",	-- 0x2f16
		"10001001",	-- 0x2f17
		"00000000",	-- 0x2f18
		"00010000",	-- 0x2f19
		"01000101",	-- 0x2f1a
		"00000101",	-- 0x2f1b
		"10000111",	-- 0x2f1c
		"00000000",	-- 0x2f1d
		"00001001",	-- 0x2f1e
		"01000000",	-- 0x2f1f
		"00000110",	-- 0x2f20
		"10000111",	-- 0x2f21
		"00000000",	-- 0x2f22
		"00000001",	-- 0x2f23
		"10001100",	-- 0x2f24
		"11001010",	-- 0x2f25
		"11111110",	-- 0x2f26
		"10111010",	-- 0x2f27
		"00000001",	-- 0x2f28
		"01011010",	-- 0x2f29
		"01000000",	-- 0x2f2a
		"00011100",	-- 0x2f2b
		"00110101",	-- 0x2f2c
		"11010000",	-- 0x2f2d
		"00011000",	-- 0x2f2e
		"00110101",	-- 0x2f2f
		"00010011",	-- 0x2f30
		"00010101",	-- 0x2f31
		"00110111",	-- 0x2f32
		"01110100",	-- 0x2f33
		"00010010",	-- 0x2f34
		"00110111",	-- 0x2f35
		"10111110",	-- 0x2f36
		"00001111",	-- 0x2f37
		"00110111",	-- 0x2f38
		"01010110",	-- 0x2f39
		"00001100",	-- 0x2f3a
		"01111001",	-- 0x2f3b
		"00000101",	-- 0x2f3c
		"01011101",	-- 0x2f3d
		"01000101",	-- 0x2f3e
		"00000111",	-- 0x2f3f
		"01111001",	-- 0x2f40
		"11000100",	-- 0x2f41
		"01010111",	-- 0x2f42
		"01000101",	-- 0x2f43
		"00000010",	-- 0x2f44
		"01110111",	-- 0x2f45
		"11011110",	-- 0x2f46
		"01100011",	-- 0x2f47
		"11011010",	-- 0x2f48
		"01001110",	-- 0x2f49
		"10110010",	-- 0x2f4a
		"00000001",	-- 0x2f4b
		"11010101",	-- 0x2f4c
		"01010010",	-- 0x2f4d
		"11111011",	-- 0x2f4e
		"00000001",	-- 0x2f4f
		"01010101",	-- 0x2f50
		"11110001",	-- 0x2f51
		"00000001",	-- 0x2f52
		"01010110",	-- 0x2f53
		"00010110",	-- 0x2f54
		"11110001",	-- 0x2f55
		"00000010",	-- 0x2f56
		"00111001",	-- 0x2f57
		"10000000",	-- 0x2f58
		"00000000",	-- 0x2f59
		"10001000",	-- 0x2f5a
		"00000000",	-- 0x2f5b
		"10000101",	-- 0x2f5c
		"01001011",	-- 0x2f5d
		"00001011",	-- 0x2f5e
		"10001001",	-- 0x2f5f
		"00000000",	-- 0x2f60
		"11100111",	-- 0x2f61
		"01000011",	-- 0x2f62
		"00000010",	-- 0x2f63
		"11001011",	-- 0x2f64
		"11100111",	-- 0x2f65
		"11001101",	-- 0x2f66
		"00000000",	-- 0x2f67
		"01000100",	-- 0x2f68
		"00000010",	-- 0x2f69
		"11001011",	-- 0x2f6a
		"00000000",	-- 0x2f6b
		"10110011",	-- 0x2f6c
		"00000001",	-- 0x2f6d
		"01010111",	-- 0x2f6e
		"11111010",	-- 0x2f6f
		"00000001",	-- 0x2f70
		"11010011",	-- 0x2f71
		"10010010",	-- 0x2f72
		"01001110",	-- 0x2f73
		"00000001",	-- 0x2f74
		"11101011",	-- 0x2f75
		"01010111",	-- 0x2f76
		"00110101",	-- 0x2f77
		"10110000",	-- 0x2f78
		"00001001",	-- 0x2f79
		"00110101",	-- 0x2f7a
		"11110110",	-- 0x2f7b
		"00000110",	-- 0x2f7c
		"00110101",	-- 0x2f7d
		"00010000",	-- 0x2f7e
		"00010101",	-- 0x2f7f
		"00110111",	-- 0x2f80
		"01111101",	-- 0x2f81
		"00000100",	-- 0x2f82
		"11001011",	-- 0x2f83
		"01000000",	-- 0x2f84
		"01000000",	-- 0x2f85
		"00001000",	-- 0x2f86
		"00110111",	-- 0x2f87
		"10111001",	-- 0x2f88
		"00001011",	-- 0x2f89
		"00110111",	-- 0x2f8a
		"01010110",	-- 0x2f8b
		"00001000",	-- 0x2f8c
		"11001011",	-- 0x2f8d
		"01000000",	-- 0x2f8e
		"10110011",	-- 0x2f8f
		"00000001",	-- 0x2f90
		"01011001",	-- 0x2f91
		"00000011",	-- 0x2f92
		"11101111",	-- 0x2f93
		"10110000",	-- 0x2f94
		"11111011",	-- 0x2f95
		"00000001",	-- 0x2f96
		"01011001",	-- 0x2f97
		"11000001",	-- 0x2f98
		"00000100",	-- 0x2f99
		"01000101",	-- 0x2f9a
		"00000101",	-- 0x2f9b
		"11111101",	-- 0x2f9c
		"00000001",	-- 0x2f9d
		"01010111",	-- 0x2f9e
		"01000011",	-- 0x2f9f
		"00000011",	-- 0x2fa0
		"11111011",	-- 0x2fa1
		"00000001",	-- 0x2fa2
		"01010111",	-- 0x2fa3
		"00110111",	-- 0x2fa4
		"00011001",	-- 0x2fa5
		"00000110",	-- 0x2fa6
		"11001101",	-- 0x2fa7
		"00101011",	-- 0x2fa8
		"01000011",	-- 0x2fa9
		"00000010",	-- 0x2faa
		"11001011",	-- 0x2fab
		"00101011",	-- 0x2fac
		"10110011",	-- 0x2fad
		"00000001",	-- 0x2fae
		"01011001",	-- 0x2faf
		"01100011",	-- 0x2fb0
		"01110101",	-- 0x2fb1
		"11001101",	-- 0x2fb2
		"01101110",	-- 0x2fb3
		"01101111",	-- 0x2fb4
		"11011011",	-- 0x2fb5
		"10100001",	-- 0x2fb6
		"01001011",	-- 0x2fb7
		"00011111",	-- 0x2fb8
		"01111001",	-- 0x2fb9
		"00111111",	-- 0x2fba
		"11000010",	-- 0x2fbb
		"01000101",	-- 0x2fbc
		"00011010",	-- 0x2fbd
		"11111010",	-- 0x2fbe
		"00000001",	-- 0x2fbf
		"10001001",	-- 0x2fc0
		"00110111",	-- 0x2fc1
		"11001100",	-- 0x2fc2
		"00000100",	-- 0x2fc3
		"01010110",	-- 0x2fc4
		"01000110",	-- 0x2fc5
		"00000001",	-- 0x2fc6
		"01010000",	-- 0x2fc7
		"00110101",	-- 0x2fc8
		"11000000",	-- 0x2fc9
		"00001110",	-- 0x2fca
		"11001100",	-- 0x2fcb
		"00000010",	-- 0x2fcc
		"01000111",	-- 0x2fcd
		"00000111",	-- 0x2fce
		"11001100",	-- 0x2fcf
		"00000110",	-- 0x2fd0
		"01000101",	-- 0x2fd1
		"00000101",	-- 0x2fd2
		"01110111",	-- 0x2fd3
		"11111011",	-- 0x2fd4
		"10001100",	-- 0x2fd5
		"01110101",	-- 0x2fd6
		"11111011",	-- 0x2fd7
		"01010010",	-- 0x2fd8
		"10110010",	-- 0x2fd9
		"00000001",	-- 0x2fda
		"10001001",	-- 0x2fdb
		"01110101",	-- 0x2fdc
		"11001100",	-- 0x2fdd
		"11011011",	-- 0x2fde
		"10100001",	-- 0x2fdf
		"00110111",	-- 0x2fe0
		"11100000",	-- 0x2fe1
		"00011110",	-- 0x2fe2
		"00110111",	-- 0x2fe3
		"11000000",	-- 0x2fe4
		"00100010",	-- 0x2fe5
		"01011001",	-- 0x2fe6
		"01001011",	-- 0x2fe7
		"00110011",	-- 0x2fe8
		"01011010",	-- 0x2fe9
		"01010111",	-- 0x2fea
		"11000010",	-- 0x2feb
		"00001111",	-- 0x2fec
		"11001100",	-- 0x2fed
		"00000101",	-- 0x2fee
		"01000101",	-- 0x2fef
		"00101011",	-- 0x2ff0
		"11000011",	-- 0x2ff1
		"11110000",	-- 0x2ff2
		"11000001",	-- 0x2ff3
		"00010000",	-- 0x2ff4
		"01011010",	-- 0x2ff5
		"11001101",	-- 0x2ff6
		"00100000",	-- 0x2ff7
		"01000111",	-- 0x2ff8
		"00010111",	-- 0x2ff9
		"11001101",	-- 0x2ffa
		"01000000",	-- 0x2ffb
		"01000110",	-- 0x2ffc
		"00011110",	-- 0x2ffd
		"01010010",	-- 0x2ffe
		"01000000",	-- 0x2fff
		"00010000",	-- 0x3000
		"01010010",	-- 0x3001
		"11001101",	-- 0x3002
		"00110101",	-- 0x3003
		"01000111",	-- 0x3004
		"00010101",	-- 0x3005
		"01000000",	-- 0x3006
		"00000110",	-- 0x3007
		"11001010",	-- 0x3008
		"00100000",	-- 0x3009
		"11001101",	-- 0x300a
		"00010101",	-- 0x300b
		"01000111",	-- 0x300c
		"00001101",	-- 0x300d
		"01011001",	-- 0x300e
		"01001011",	-- 0x300f
		"00001010",	-- 0x3010
		"00110111",	-- 0x3011
		"01010000",	-- 0x3012
		"00000111",	-- 0x3013
		"00110101",	-- 0x3014
		"00010110",	-- 0x3015
		"00000100",	-- 0x3016
		"01110111",	-- 0x3017
		"01111000",	-- 0x3018
		"01110111",	-- 0x3019
		"00111011",	-- 0x301a
		"01011011",	-- 0x301b
		"10010011",	-- 0x301c
		"10100001",	-- 0x301d
		"01000000",	-- 0x301e
		"00101111",	-- 0x301f
		"10000110",	-- 0x3020
		"01010101",	-- 0x3021
		"00000000",	-- 0x3022
		"10001111",	-- 0x3023
		"00000000",	-- 0x3024
		"11110000",	-- 0x3025
		"10001010",	-- 0x3026
		"10001010",	-- 0x3027
		"10001010",	-- 0x3028
		"10000110",	-- 0x3029
		"11111111",	-- 0x302a
		"11111111",	-- 0x302b
		"10011010",	-- 0x302c
		"11110110",	-- 0x302d
		"10010010",	-- 0x302e
		"10100001",	-- 0x302f
		"10010010",	-- 0x3030
		"10100010",	-- 0x3031
		"01100011",	-- 0x3032
		"00110111",	-- 0x3033
		"00011001",	-- 0x3034
		"00010001",	-- 0x3035
		"01110001",	-- 0x3036
		"11110100",	-- 0x3037
		"01000110",	-- 0x3038
		"00010100",	-- 0x3039
		"01111001",	-- 0x303a
		"00001100",	-- 0x303b
		"10101110",	-- 0x303c
		"01000101",	-- 0x303d
		"00001111",	-- 0x303e
		"11001010",	-- 0x303f
		"11111111",	-- 0x3040
		"10010010",	-- 0x3041
		"10100001",	-- 0x3042
		"10010010",	-- 0x3043
		"10100010",	-- 0x3044
		"01000000",	-- 0x3045
		"00000111",	-- 0x3046
		"00110111",	-- 0x3047
		"11110100",	-- 0x3048
		"00000100",	-- 0x3049
		"01110101",	-- 0x304a
		"11110100",	-- 0x304b
		"01110010",	-- 0x304c
		"10101110",	-- 0x304d
		"01100011",	-- 0x304e
		"00000001",	-- 0x304f
		"11110100",	-- 0x3050
		"01101111",	-- 0x3051
		"01110101",	-- 0x3052
		"01110010",	-- 0x3053
		"01110111",	-- 0x3054
		"00101101",	-- 0x3055
		"01111111",	-- 0x3056
		"01111110",	-- 0x3057
		"01110011",	-- 0x3058
		"00000001",	-- 0x3059
		"11001101",	-- 0x305a
		"00110101",	-- 0x305b
		"00000001",	-- 0x305c
		"11011101",	-- 0x305d
		"00101010",	-- 0x305e
		"10011110",	-- 0x305f
		"00011000",	-- 0x3060
		"00001010",	-- 0x3061
		"00000001",	-- 0x3062
		"00000101",	-- 0x3063
		"01010010",	-- 0x3064
		"11011011",	-- 0x3065
		"10100001",	-- 0x3066
		"01001010",	-- 0x3067
		"00000010",	-- 0x3068
		"11001010",	-- 0x3069
		"00001000",	-- 0x306a
		"01111010",	-- 0x306b
		"11000111",	-- 0x306c
		"01111011",	-- 0x306d
		"10100010",	-- 0x306e
		"01011001",	-- 0x306f
		"01001011",	-- 0x3070
		"00011100",	-- 0x3071
		"11011011",	-- 0x3072
		"10100010",	-- 0x3073
		"11000011",	-- 0x3074
		"00000111",	-- 0x3075
		"11001111",	-- 0x3076
		"00000001",	-- 0x3077
		"01000110",	-- 0x3078
		"00011111",	-- 0x3079
		"10001111",	-- 0x307a
		"00000000",	-- 0x307b
		"11110000",	-- 0x307c
		"00001111",	-- 0x307d
		"11001100",	-- 0x307e
		"00001000",	-- 0x307f
		"01000100",	-- 0x3080
		"00001000",	-- 0x3081
		"00111100",	-- 0x3082
		"10111000",	-- 0x3083
		"00000001",	-- 0x3084
		"00000111",	-- 0x3085
		"11001100",	-- 0x3086
		"01010101",	-- 0x3087
		"01000101",	-- 0x3088
		"00000011",	-- 0x3089
		"10000110",	-- 0x308a
		"01010101",	-- 0x308b
		"00000000",	-- 0x308c
		"10001010",	-- 0x308d
		"00001010",	-- 0x308e
		"00000001",	-- 0x308f
		"00000111",	-- 0x3090
		"10010110",	-- 0x3091
		"11110000",	-- 0x3092
		"10010111",	-- 0x3093
		"11110010",	-- 0x3094
		"10010111",	-- 0x3095
		"11110100",	-- 0x3096
		"10011010",	-- 0x3097
		"11110110",	-- 0x3098
		"11011011",	-- 0x3099
		"10100010",	-- 0x309a
		"01001010",	-- 0x309b
		"00000011",	-- 0x309c
		"00000011",	-- 0x309d
		"11110010",	-- 0x309e
		"01101111",	-- 0x309f
		"11000011",	-- 0x30a0
		"00000111",	-- 0x30a1
		"01101101",	-- 0x30a2
		"01000110",	-- 0x30a3
		"00000010",	-- 0x30a4
		"01110101",	-- 0x30a5
		"00110001",	-- 0x30a6
		"11001101",	-- 0x30a7
		"00000100",	-- 0x30a8
		"01000110",	-- 0x30a9
		"00110100",	-- 0x30aa
		"00110101",	-- 0x30ab
		"01010101",	-- 0x30ac
		"00110001",	-- 0x30ad
		"01111001",	-- 0x30ae
		"00111100",	-- 0x30af
		"01011011",	-- 0x30b0
		"01000100",	-- 0x30b1
		"00101100",	-- 0x30b2
		"11001010",	-- 0x30b3
		"00000010",	-- 0x30b4
		"11001011",	-- 0x30b5
		"01010110",	-- 0x30b6
		"10111000",	-- 0x30b7
		"00000001",	-- 0x30b8
		"01110101",	-- 0x30b9
		"00000100",	-- 0x30ba
		"10010010",	-- 0x30bb
		"10100100",	-- 0x30bc
		"10011110",	-- 0x30bd
		"11110100",	-- 0x30be
		"00000001",	-- 0x30bf
		"11000101",	-- 0x30c0
		"01011010",	-- 0x30c1
		"01111001",	-- 0x30c2
		"00000000",	-- 0x30c3
		"10100100",	-- 0x30c4
		"01000111",	-- 0x30c5
		"00000010",	-- 0x30c6
		"10010111",	-- 0x30c7
		"11110100",	-- 0x30c8
		"10001000",	-- 0x30c9
		"00000000",	-- 0x30ca
		"00110101",	-- 0x30cb
		"10110111",	-- 0x30cc
		"00000001",	-- 0x30cd
		"00000111",	-- 0x30ce
		"10111000",	-- 0x30cf
		"00000001",	-- 0x30d0
		"01110011",	-- 0x30d1
		"00111110",	-- 0x30d2
		"00000101",	-- 0x30d3
		"10011001",	-- 0x30d4
		"00001000",	-- 0x30d5
		"01001010",	-- 0x30d6
		"00000110",	-- 0x30d7
		"00110111",	-- 0x30d8
		"00010101",	-- 0x30d9
		"00000011",	-- 0x30da
		"00000001",	-- 0x30db
		"11110010",	-- 0x30dc
		"00101001",	-- 0x30dd
		"00000111",	-- 0x30de
		"01111101",	-- 0x30df
		"00110111",	-- 0x30e0
		"01010101",	-- 0x30e1
		"00101000",	-- 0x30e2
		"11001101",	-- 0x30e3
		"00000011",	-- 0x30e4
		"01000110",	-- 0x30e5
		"00000010",	-- 0x30e6
		"01110101",	-- 0x30e7
		"10010101",	-- 0x30e8
		"00110101",	-- 0x30e9
		"10010101",	-- 0x30ea
		"00011100",	-- 0x30eb
		"11001010",	-- 0x30ec
		"00101011",	-- 0x30ed
		"10110010",	-- 0x30ee
		"00000001",	-- 0x30ef
		"01101111",	-- 0x30f0
		"11001010",	-- 0x30f1
		"01001011",	-- 0x30f2
		"10110010",	-- 0x30f3
		"00000010",	-- 0x30f4
		"00011000",	-- 0x30f5
		"01011001",	-- 0x30f6
		"01000110",	-- 0x30f7
		"00000101",	-- 0x30f8
		"00000101",	-- 0x30f9
		"01110101",	-- 0x30fa
		"00000110",	-- 0x30fb
		"01000000",	-- 0x30fc
		"00000111",	-- 0x30fd
		"11001101",	-- 0x30fe
		"00000101",	-- 0x30ff
		"01000110",	-- 0x3100
		"00000110",	-- 0x3101
		"00000101",	-- 0x3102
		"01110111",	-- 0x3103
		"00000110",	-- 0x3104
		"00000001",	-- 0x3105
		"11110010",	-- 0x3106
		"01011010",	-- 0x3107
		"00000011",	-- 0x3108
		"11110010",	-- 0x3109
		"01101111",	-- 0x310a
		"00111111",	-- 0x310b
		"11001101",	-- 0x310c
		"00000001",	-- 0x310d
		"01000111",	-- 0x310e
		"00000111",	-- 0x310f
		"11001101",	-- 0x3110
		"00000011",	-- 0x3111
		"01000111",	-- 0x3112
		"00001010",	-- 0x3113
		"00000011",	-- 0x3114
		"11110001",	-- 0x3115
		"11100111",	-- 0x3116
		"11111011",	-- 0x3117
		"00000001",	-- 0x3118
		"01011001",	-- 0x3119
		"01110101",	-- 0x311a
		"10110101",	-- 0x311b
		"01000000",	-- 0x311c
		"00000011",	-- 0x311d
		"11111011",	-- 0x311e
		"00000001",	-- 0x311f
		"01101111",	-- 0x3120
		"01110101",	-- 0x3121
		"10010101",	-- 0x3122
		"00110101",	-- 0x3123
		"11110110",	-- 0x3124
		"00010001",	-- 0x3125
		"00110101",	-- 0x3126
		"00010000",	-- 0x3127
		"00011001",	-- 0x3128
		"00110101",	-- 0x3129
		"01111101",	-- 0x312a
		"00001011",	-- 0x312b
		"00110111",	-- 0x312c
		"01010110",	-- 0x312d
		"00010011",	-- 0x312e
		"00110111",	-- 0x312f
		"10111001",	-- 0x3130
		"00010000",	-- 0x3131
		"10000110",	-- 0x3132
		"00000000",	-- 0x3133
		"10000000",	-- 0x3134
		"01000000",	-- 0x3135
		"00000011",	-- 0x3136
		"10000110",	-- 0x3137
		"00000000",	-- 0x3138
		"01010110",	-- 0x3139
		"00111110",	-- 0x313a
		"00000100",	-- 0x313b
		"10110011",	-- 0x313c
		"00000001",	-- 0x313d
		"01101111",	-- 0x313e
		"00111100",	-- 0x313f
		"01000000",	-- 0x3140
		"01000111",	-- 0x3141
		"11111101",	-- 0x3142
		"00000001",	-- 0x3143
		"01011101",	-- 0x3144
		"01000101",	-- 0x3145
		"00000011",	-- 0x3146
		"11111011",	-- 0x3147
		"00000001",	-- 0x3148
		"01011101",	-- 0x3149
		"01010010",	-- 0x314a
		"00000110",	-- 0x314b
		"10011010",	-- 0x314c
		"10100100",	-- 0x314d
		"01010010",	-- 0x314e
		"11111011",	-- 0x314f
		"00000001",	-- 0x3150
		"01010111",	-- 0x3151
		"00000110",	-- 0x3152
		"11110101",	-- 0x3153
		"00000010",	-- 0x3154
		"00011011",	-- 0x3155
		"10000100",	-- 0x3156
		"00000000",	-- 0x3157
		"01000100",	-- 0x3158
		"00000010",	-- 0x3159
		"01010010",	-- 0x315a
		"01010011",	-- 0x315b
		"10011001",	-- 0x315c
		"10100100",	-- 0x315d
		"01000101",	-- 0x315e
		"00000010",	-- 0x315f
		"10010110",	-- 0x3160
		"10100100",	-- 0x3161
		"10111001",	-- 0x3162
		"00000001",	-- 0x3163
		"01011010",	-- 0x3164
		"01000101",	-- 0x3165
		"00000011",	-- 0x3166
		"10110110",	-- 0x3167
		"00000001",	-- 0x3168
		"01011010",	-- 0x3169
		"00111110",	-- 0x316a
		"00000100",	-- 0x316b
		"10110011",	-- 0x316c
		"00000001",	-- 0x316d
		"01101111",	-- 0x316e
		"11111010",	-- 0x316f
		"00000001",	-- 0x3170
		"01011000",	-- 0x3171
		"00001100",	-- 0x3172
		"00111100",	-- 0x3173
		"10001000",	-- 0x3174
		"00000000",	-- 0x3175
		"01010101",	-- 0x3176
		"01000100",	-- 0x3177
		"00000010",	-- 0x3178
		"01010010",	-- 0x3179
		"01010011",	-- 0x317a
		"00111110",	-- 0x317b
		"11111010",	-- 0x317c
		"00000010",	-- 0x317d
		"01000110",	-- 0x317e
		"01111001",	-- 0x317f
		"00110000",	-- 0x3180
		"10100010",	-- 0x3181
		"01000100",	-- 0x3182
		"00000011",	-- 0x3183
		"11111010",	-- 0x3184
		"00000010",	-- 0x3185
		"01000111",	-- 0x3186
		"00001100",	-- 0x3187
		"00111100",	-- 0x3188
		"10001001",	-- 0x3189
		"00000001",	-- 0x318a
		"11001101",	-- 0x318b
		"01000011",	-- 0x318c
		"00000011",	-- 0x318d
		"10000110",	-- 0x318e
		"00000001",	-- 0x318f
		"11001101",	-- 0x3190
		"00111110",	-- 0x3191
		"00000100",	-- 0x3192
		"00010001",	-- 0x3193
		"11000001",	-- 0x3194
		"00110101",	-- 0x3195
		"10110011",	-- 0x3196
		"00000010",	-- 0x3197
		"00011000",	-- 0x3198
		"00111100",	-- 0x3199
		"10001000",	-- 0x319a
		"00000000",	-- 0x319b
		"00000111",	-- 0x319c
		"01000100",	-- 0x319d
		"00000010",	-- 0x319e
		"01010010",	-- 0x319f
		"01010011",	-- 0x31a0
		"10111010",	-- 0x31a1
		"00000001",	-- 0x31a2
		"01110101",	-- 0x31a3
		"00111101",	-- 0x31a4
		"11001010",	-- 0x31a5
		"00000110",	-- 0x31a6
		"00001001",	-- 0x31a7
		"11001011",	-- 0x31a8
		"01010110",	-- 0x31a9
		"10111000",	-- 0x31aa
		"00000001",	-- 0x31ab
		"01110101",	-- 0x31ac
		"00111110",	-- 0x31ad
		"11011010",	-- 0x31ae
		"01011001",	-- 0x31af
		"10000001",	-- 0x31b0
		"11101001",	-- 0x31b1
		"10010010",	-- 0x31b2
		"10100100",	-- 0x31b3
		"00111100",	-- 0x31b4
		"00010001",	-- 0x31b5
		"11011101",	-- 0x31b6
		"10100100",	-- 0x31b7
		"01000100",	-- 0x31b8
		"00001001",	-- 0x31b9
		"01010000",	-- 0x31ba
		"01001010",	-- 0x31bb
		"00000100",	-- 0x31bc
		"01010010",	-- 0x31bd
		"11011011",	-- 0x31be
		"10100100",	-- 0x31bf
		"10001100",	-- 0x31c0
		"11000001",	-- 0x31c1
		"10000000",	-- 0x31c2
		"01010110",	-- 0x31c3
		"10111010",	-- 0x31c4
		"00000001",	-- 0x31c5
		"01101011",	-- 0x31c6
		"00111100",	-- 0x31c7
		"10010011",	-- 0x31c8
		"10100100",	-- 0x31c9
		"01011011",	-- 0x31ca
		"01010010",	-- 0x31cb
		"10000101",	-- 0x31cc
		"00000110",	-- 0x31cd
		"01111011",	-- 0x31ce
		"10100100",	-- 0x31cf
		"10000101",	-- 0x31d0
		"00000110",	-- 0x31d1
		"01011010",	-- 0x31d2
		"00000001",	-- 0x31d3
		"11110010",	-- 0x31d4
		"01100011",	-- 0x31d5
		"01111001",	-- 0x31d6
		"00000000",	-- 0x31d7
		"10100100",	-- 0x31d8
		"01000111",	-- 0x31d9
		"00000010",	-- 0x31da
		"10010111",	-- 0x31db
		"11110110",	-- 0x31dc
		"10001000",	-- 0x31dd
		"00000000",	-- 0x31de
		"00110101",	-- 0x31df
		"10110111",	-- 0x31e0
		"00000001",	-- 0x31e1
		"00000101",	-- 0x31e2
		"01100001",	-- 0x31e3
		"00100100",	-- 0x31e4
		"01110111",	-- 0x31e5
		"00010101",	-- 0x31e6
		"10110110",	-- 0x31e7
		"00000001",	-- 0x31e8
		"01101011",	-- 0x31e9
		"01010000",	-- 0x31ea
		"10110010",	-- 0x31eb
		"00000001",	-- 0x31ec
		"01101011",	-- 0x31ed
		"01000110",	-- 0x31ee
		"01111111",	-- 0x31ef
		"01011010",	-- 0x31f0
		"01100001",	-- 0x31f1
		"01110000",	-- 0x31f2
		"10010011",	-- 0x31f3
		"10100100",	-- 0x31f4
		"01011011",	-- 0x31f5
		"01010010",	-- 0x31f6
		"10000101",	-- 0x31f7
		"00000011",	-- 0x31f8
		"01111011",	-- 0x31f9
		"10100100",	-- 0x31fa
		"10000101",	-- 0x31fb
		"00000011",	-- 0x31fc
		"11011010",	-- 0x31fd
		"10100100",	-- 0x31fe
		"10001000",	-- 0x31ff
		"00000000",	-- 0x3200
		"00110101",	-- 0x3201
		"10110111",	-- 0x3202
		"00000001",	-- 0x3203
		"00000101",	-- 0x3204
		"01100001",	-- 0x3205
		"00111001",	-- 0x3206
		"01000000",	-- 0x3207
		"01100110",	-- 0x3208
		"10111000",	-- 0x3209
		"00000001",	-- 0x320a
		"01110011",	-- 0x320b
		"00111110",	-- 0x320c
		"01111001",	-- 0x320d
		"00011101",	-- 0x320e
		"11110110",	-- 0x320f
		"01000100",	-- 0x3210
		"00010111",	-- 0x3211
		"10111000",	-- 0x3212
		"00000001",	-- 0x3213
		"01110000",	-- 0x3214
		"01001011",	-- 0x3215
		"00001001",	-- 0x3216
		"00000100",	-- 0x3217
		"01011000",	-- 0x3218
		"01000110",	-- 0x3219
		"00001110",	-- 0x321a
		"11111101",	-- 0x321b
		"00000001",	-- 0x321c
		"01110010",	-- 0x321d
		"01000100",	-- 0x321e
		"00001001",	-- 0x321f
		"01010010",	-- 0x3220
		"11111011",	-- 0x3221
		"00000001",	-- 0x3222
		"01110010",	-- 0x3223
		"00000110",	-- 0x3224
		"10110111",	-- 0x3225
		"00000001",	-- 0x3226
		"01110000",	-- 0x3227
		"00111110",	-- 0x3228
		"00001010",	-- 0x3229
		"00000001",	-- 0x322a
		"01101001",	-- 0x322b
		"00000101",	-- 0x322c
		"00110111",	-- 0x322d
		"00000110",	-- 0x322e
		"00001100",	-- 0x322f
		"10010110",	-- 0x3230
		"00000100",	-- 0x3231
		"10000111",	-- 0x3232
		"00000000",	-- 0x3233
		"00000100",	-- 0x3234
		"10011001",	-- 0x3235
		"00001000",	-- 0x3236
		"01001010",	-- 0x3237
		"00101000",	-- 0x3238
		"01010110",	-- 0x3239
		"10011010",	-- 0x323a
		"00001000",	-- 0x323b
		"01110111",	-- 0x323c
		"00000110",	-- 0x323d
		"01000000",	-- 0x323e
		"00010000",	-- 0x323f
		"10111010",	-- 0x3240
		"00000001",	-- 0x3241
		"01101001",	-- 0x3242
		"00000101",	-- 0x3243
		"00110101",	-- 0x3244
		"01110101",	-- 0x3245
		"00000100",	-- 0x3246
		"01110111",	-- 0x3247
		"10110101",	-- 0x3248
		"01000000",	-- 0x3249
		"00010110",	-- 0x324a
		"00000101",	-- 0x324b
		"01110101",	-- 0x324c
		"00000110",	-- 0x324d
		"01110101",	-- 0x324e
		"00110101",	-- 0x324f
		"10110110",	-- 0x3250
		"00000001",	-- 0x3251
		"01101001",	-- 0x3252
		"10001000",	-- 0x3253
		"00000000",	-- 0x3254
		"00000100",	-- 0x3255
		"10011001",	-- 0x3256
		"00000100",	-- 0x3257
		"01001010",	-- 0x3258
		"00000010",	-- 0x3259
		"10010110",	-- 0x325a
		"00000100",	-- 0x325b
		"10000111",	-- 0x325c
		"00000000",	-- 0x325d
		"00000100",	-- 0x325e
		"10011010",	-- 0x325f
		"00001000",	-- 0x3260
		"00000111",	-- 0x3261
		"01100011",	-- 0x3262
		"00111111",	-- 0x3263
		"10010001",	-- 0x3264
		"11110110",	-- 0x3265
		"00111110",	-- 0x3266
		"00111101",	-- 0x3267
		"10010001",	-- 0x3268
		"11110111",	-- 0x3269
		"10000000",	-- 0x326a
		"00000000",	-- 0x326b
		"00001100",	-- 0x326c
		"00111100",	-- 0x326d
		"01100011",	-- 0x326e
		"11011010",	-- 0x326f
		"10100010",	-- 0x3270
		"01001010",	-- 0x3271
		"00000011",	-- 0x3272
		"00000011",	-- 0x3273
		"11110011",	-- 0x3274
		"10101111",	-- 0x3275
		"10110110",	-- 0x3276
		"00000001",	-- 0x3277
		"00001010",	-- 0x3278
		"00110101",	-- 0x3279
		"00010110",	-- 0x327a
		"00100001",	-- 0x327b
		"00110101",	-- 0x327c
		"10110100",	-- 0x327d
		"01010011",	-- 0x327e
		"01111001",	-- 0x327f
		"00011000",	-- 0x3280
		"01011011",	-- 0x3281
		"01000100",	-- 0x3282
		"00000101",	-- 0x3283
		"01111001",	-- 0x3284
		"00011111",	-- 0x3285
		"11010000",	-- 0x3286
		"01000101",	-- 0x3287
		"00010100",	-- 0x3288
		"01111001",	-- 0x3289
		"00010001",	-- 0x328a
		"10100010",	-- 0x328b
		"01000110",	-- 0x328c
		"00001111",	-- 0x328d
		"00000100",	-- 0x328e
		"01110111",	-- 0x328f
		"10110100",	-- 0x3290
		"10001110",	-- 0x3291
		"11110011",	-- 0x3292
		"01101001",	-- 0x3293
		"00000001",	-- 0x3294
		"11110011",	-- 0x3295
		"11100111",	-- 0x3296
		"00011100",	-- 0x3297
		"00000001",	-- 0x3298
		"11110011",	-- 0x3299
		"11100111",	-- 0x329a
		"01000000",	-- 0x329b
		"00101001",	-- 0x329c
		"01110101",	-- 0x329d
		"10110100",	-- 0x329e
		"10001110",	-- 0x329f
		"11110011",	-- 0x32a0
		"01101001",	-- 0x32a1
		"01111001",	-- 0x32a2
		"00010010",	-- 0x32a3
		"10100010",	-- 0x32a4
		"01000111",	-- 0x32a5
		"00010011",	-- 0x32a6
		"01111001",	-- 0x32a7
		"00110010",	-- 0x32a8
		"10100010",	-- 0x32a9
		"01000111",	-- 0x32aa
		"00001110",	-- 0x32ab
		"00011100",	-- 0x32ac
		"01111001",	-- 0x32ad
		"00000010",	-- 0x32ae
		"10100010",	-- 0x32af
		"01000111",	-- 0x32b0
		"00001000",	-- 0x32b1
		"01111001",	-- 0x32b2
		"00100010",	-- 0x32b3
		"10100010",	-- 0x32b4
		"01000111",	-- 0x32b5
		"00000011",	-- 0x32b6
		"00000011",	-- 0x32b7
		"11110011",	-- 0x32b8
		"01000101",	-- 0x32b9
		"00110111",	-- 0x32ba
		"11110101",	-- 0x32bb
		"00000001",	-- 0x32bc
		"00000100",	-- 0x32bd
		"00000001",	-- 0x32be
		"11110011",	-- 0x32bf
		"11100111",	-- 0x32c0
		"00011100",	-- 0x32c1
		"00011100",	-- 0x32c2
		"00000001",	-- 0x32c3
		"11110011",	-- 0x32c4
		"11100111",	-- 0x32c5
		"11001010",	-- 0x32c6
		"00000010",	-- 0x32c7
		"10110010",	-- 0x32c8
		"00000001",	-- 0x32c9
		"01001011",	-- 0x32ca
		"11001010",	-- 0x32cb
		"00010000",	-- 0x32cc
		"10110010",	-- 0x32cd
		"00000001",	-- 0x32ce
		"01001101",	-- 0x32cf
		"01000000",	-- 0x32d0
		"01010100",	-- 0x32d1
		"11111011",	-- 0x32d2
		"00000001",	-- 0x32d3
		"01001110",	-- 0x32d4
		"01011010",	-- 0x32d5
		"11001101",	-- 0x32d6
		"00110101",	-- 0x32d7
		"01000010",	-- 0x32d8
		"11101100",	-- 0x32d9
		"11000011",	-- 0x32da
		"00001111",	-- 0x32db
		"11001101",	-- 0x32dc
		"00000101",	-- 0x32dd
		"01000010",	-- 0x32de
		"11100110",	-- 0x32df
		"11011100",	-- 0x32e0
		"10100010",	-- 0x32e1
		"01000110",	-- 0x32e2
		"01100001",	-- 0x32e3
		"11111011",	-- 0x32e4
		"00000001",	-- 0x32e5
		"01001011",	-- 0x32e6
		"11000011",	-- 0x32e7
		"00000011",	-- 0x32e8
		"10001110",	-- 0x32e9
		"11110011",	-- 0x32ea
		"01101001",	-- 0x32eb
		"00001110",	-- 0x32ec
		"10001111",	-- 0x32ed
		"00000001",	-- 0x32ee
		"00001010",	-- 0x32ef
		"00001111",	-- 0x32f0
		"00001111",	-- 0x32f1
		"10100110",	-- 0x32f2
		"10000000",	-- 0x32f3
		"00000001",	-- 0x32f4
		"11110011",	-- 0x32f5
		"11100111",	-- 0x32f6
		"11111010",	-- 0x32f7
		"00000001",	-- 0x32f8
		"01001011",	-- 0x32f9
		"01010110",	-- 0x32fa
		"11000010",	-- 0x32fb
		"00000011",	-- 0x32fc
		"10110010",	-- 0x32fd
		"00000001",	-- 0x32fe
		"01001011",	-- 0x32ff
		"10110110",	-- 0x3300
		"00000001",	-- 0x3301
		"01001100",	-- 0x3302
		"00001001",	-- 0x3303
		"01000101",	-- 0x3304
		"00001000",	-- 0x3305
		"11001100",	-- 0x3306
		"00000101",	-- 0x3307
		"01000011",	-- 0x3308
		"00011000",	-- 0x3309
		"11001010",	-- 0x330a
		"00000101",	-- 0x330b
		"01000000",	-- 0x330c
		"00010100",	-- 0x330d
		"11001100",	-- 0x330e
		"11111101",	-- 0x330f
		"01000100",	-- 0x3310
		"00001010",	-- 0x3311
		"01101101",	-- 0x3312
		"11111011",	-- 0x3313
		"00000001",	-- 0x3314
		"01001011",	-- 0x3315
		"00010001",	-- 0x3316
		"01111101",	-- 0x3317
		"01000101",	-- 0x3318
		"00000010",	-- 0x3319
		"01110101",	-- 0x331a
		"01110001",	-- 0x331b
		"11001100",	-- 0x331c
		"11111011",	-- 0x331d
		"01000100",	-- 0x331e
		"00000010",	-- 0x331f
		"11001010",	-- 0x3320
		"11111011",	-- 0x3321
		"00001000",	-- 0x3322
		"10110010",	-- 0x3323
		"00000001",	-- 0x3324
		"01001101",	-- 0x3325
		"11111010",	-- 0x3326
		"00000001",	-- 0x3327
		"01001011",	-- 0x3328
		"10000001",	-- 0x3329
		"00000110",	-- 0x332a
		"11110001",	-- 0x332b
		"00000001",	-- 0x332c
		"01001101",	-- 0x332d
		"11000101",	-- 0x332e
		"00001100",	-- 0x332f
		"01000100",	-- 0x3330
		"00000010",	-- 0x3331
		"11000001",	-- 0x3332
		"00011000",	-- 0x3333
		"11001101",	-- 0x3334
		"00011000",	-- 0x3335
		"01000101",	-- 0x3336
		"00000010",	-- 0x3337
		"11000101",	-- 0x3338
		"00011000",	-- 0x3339
		"01010010",	-- 0x333a
		"10000101",	-- 0x333b
		"00000110",	-- 0x333c
		"00010011",	-- 0x333d
		"00010011",	-- 0x333e
		"00010011",	-- 0x333f
		"00010011",	-- 0x3340
		"00001000",	-- 0x3341
		"10110010",	-- 0x3342
		"00000001",	-- 0x3343
		"01001110",	-- 0x3344
		"00110111",	-- 0x3345
		"10110100",	-- 0x3346
		"00011101",	-- 0x3347
		"11111010",	-- 0x3348
		"00000001",	-- 0x3349
		"01001110",	-- 0x334a
		"01011011",	-- 0x334b
		"11000010",	-- 0x334c
		"00000111",	-- 0x334d
		"11000011",	-- 0x334e
		"00110000",	-- 0x334f
		"11000100",	-- 0x3350
		"00000011",	-- 0x3351
		"01000100",	-- 0x3352
		"00000110",	-- 0x3353
		"11000101",	-- 0x3354
		"00010000",	-- 0x3355
		"11000011",	-- 0x3356
		"00110000",	-- 0x3357
		"11000000",	-- 0x3358
		"00000110",	-- 0x3359
		"00001000",	-- 0x335a
		"11011100",	-- 0x335b
		"10100010",	-- 0x335c
		"01000110",	-- 0x335d
		"00001000",	-- 0x335e
		"11111010",	-- 0x335f
		"00000001",	-- 0x3360
		"01001011",	-- 0x3361
		"00010000",	-- 0x3362
		"01000101",	-- 0x3363
		"00000010",	-- 0x3364
		"01110101",	-- 0x3365
		"01110001",	-- 0x3366
		"01000000",	-- 0x3367
		"01000110",	-- 0x3368
		"00010000",	-- 0x3369
		"01000000",	-- 0x336a
		"10000000",	-- 0x336b
		"00100000",	-- 0x336c
		"11101111",	-- 0x336d
		"10111111",	-- 0x336e
		"01111111",	-- 0x336f
		"11011111",	-- 0x3370
		"00111000",	-- 0x3371
		"00111100",	-- 0x3372
		"00111110",	-- 0x3373
		"00111010",	-- 0x3374
		"10110110",	-- 0x3375
		"00000001",	-- 0x3376
		"00001010",	-- 0x3377
		"10000111",	-- 0x3378
		"00000101",	-- 0x3379
		"10010001",	-- 0x337a
		"00010100",	-- 0x337b
		"00010101",	-- 0x337c
		"00000001",	-- 0x337d
		"11000100",	-- 0x337e
		"11001100",	-- 0x337f
		"00111110",	-- 0x3380
		"10010110",	-- 0x3381
		"01011001",	-- 0x3382
		"00000001",	-- 0x3383
		"11000100",	-- 0x3384
		"11001100",	-- 0x3385
		"00000001",	-- 0x3386
		"11000101",	-- 0x3387
		"00000111",	-- 0x3388
		"10000101",	-- 0x3389
		"00110001",	-- 0x338a
		"10001111",	-- 0x338b
		"11000010",	-- 0x338c
		"01100011",	-- 0x338d
		"00110101",	-- 0x338e
		"01010110",	-- 0x338f
		"00000010",	-- 0x3390
		"00011101",	-- 0x3391
		"00011101",	-- 0x3392
		"01111001",	-- 0x3393
		"10110011",	-- 0x3394
		"01010111",	-- 0x3395
		"01000101",	-- 0x3396
		"00000001",	-- 0x3397
		"00011101",	-- 0x3398
		"11101010",	-- 0x3399
		"10000000",	-- 0x339a
		"10110010",	-- 0x339b
		"00000001",	-- 0x339c
		"00001001",	-- 0x339d
		"11100001",	-- 0x339e
		"10000000",	-- 0x339f
		"11001101",	-- 0x33a0
		"00011010",	-- 0x33a1
		"01000011",	-- 0x33a2
		"00000010",	-- 0x33a3
		"11001011",	-- 0x33a4
		"00011010",	-- 0x33a5
		"11000101",	-- 0x33a6
		"00011000",	-- 0x33a7
		"01010101",	-- 0x33a8
		"11000001",	-- 0x33a9
		"00001010",	-- 0x33aa
		"10110011",	-- 0x33ab
		"00000001",	-- 0x33ac
		"01001100",	-- 0x33ad
		"01100011",	-- 0x33ae
		"00000001",	-- 0x33af
		"11110101",	-- 0x33b0
		"00101010",	-- 0x33b1
		"11011010",	-- 0x33b2
		"10100010",	-- 0x33b3
		"11001100",	-- 0x33b4
		"00000000",	-- 0x33b5
		"01000111",	-- 0x33b6
		"00000100",	-- 0x33b7
		"11001100",	-- 0x33b8
		"00100000",	-- 0x33b9
		"01000110",	-- 0x33ba
		"00000010",	-- 0x33bb
		"01110101",	-- 0x33bc
		"01010001",	-- 0x33bd
		"11000010",	-- 0x33be
		"00000111",	-- 0x33bf
		"01000110",	-- 0x33c0
		"00001010",	-- 0x33c1
		"01110101",	-- 0x33c2
		"00010001",	-- 0x33c3
		"01110101",	-- 0x33c4
		"00110100",	-- 0x33c5
		"00000001",	-- 0x33c6
		"11101101",	-- 0x33c7
		"11001011",	-- 0x33c8
		"00000001",	-- 0x33c9
		"11001110",	-- 0x33ca
		"00101001",	-- 0x33cb
		"01100011",	-- 0x33cc
		"00000001",	-- 0x33cd
		"11110100",	-- 0x33ce
		"01100000",	-- 0x33cf
		"01000000",	-- 0x33d0
		"00000011",	-- 0x33d1
		"00000001",	-- 0x33d2
		"11110100",	-- 0x33d3
		"01011011",	-- 0x33d4
		"01000100",	-- 0x33d5
		"00000011",	-- 0x33d6
		"00000011",	-- 0x33d7
		"11110100",	-- 0x33d8
		"01011010",	-- 0x33d9
		"10001110",	-- 0x33da
		"11110011",	-- 0x33db
		"01101001",	-- 0x33dc
		"01100001",	-- 0x33dd
		"00100001",	-- 0x33de
		"00011100",	-- 0x33df
		"10001100",	-- 0x33e0
		"11110011",	-- 0x33e1
		"01101100",	-- 0x33e2
		"01000011",	-- 0x33e3
		"11111000",	-- 0x33e4
		"01000000",	-- 0x33e5
		"01110011",	-- 0x33e6
		"01100001",	-- 0x33e7
		"01110111",	-- 0x33e8
		"01000101",	-- 0x33e9
		"01101111",	-- 0x33ea
		"10001001",	-- 0x33eb
		"00000000",	-- 0x33ec
		"00001101",	-- 0x33ed
		"01000101",	-- 0x33ee
		"01101010",	-- 0x33ef
		"00111111",	-- 0x33f0
		"11111010",	-- 0x33f1
		"00000001",	-- 0x33f2
		"11011100",	-- 0x33f3
		"11000110",	-- 0x33f4
		"00000010",	-- 0x33f5
		"10110010",	-- 0x33f6
		"00000001",	-- 0x33f7
		"11011100",	-- 0x33f8
		"00111101",	-- 0x33f9
		"01000000",	-- 0x33fa
		"00001001",	-- 0x33fb
		"01100001",	-- 0x33fc
		"01011101",	-- 0x33fd
		"01000101",	-- 0x33fe
		"01011010",	-- 0x33ff
		"10001001",	-- 0x3400
		"00000000",	-- 0x3401
		"00001101",	-- 0x3402
		"01000101",	-- 0x3403
		"01010101",	-- 0x3404
		"01101000",	-- 0x3405
		"01010010",	-- 0x3406
		"11101011",	-- 0x3407
		"00001000",	-- 0x3408
		"00111111",	-- 0x3409
		"00000101",	-- 0x340a
		"11011010",	-- 0x340b
		"00100101",	-- 0x340c
		"11101110",	-- 0x340d
		"00000000",	-- 0x340e
		"01000110",	-- 0x340f
		"00001000",	-- 0x3410
		"01111000",	-- 0x3411
		"01101000",	-- 0x3412
		"10110111",	-- 0x3413
		"00000001",	-- 0x3414
		"00011010",	-- 0x3415
		"01101110",	-- 0x3416
		"01000000",	-- 0x3417
		"00001110",	-- 0x3418
		"10100110",	-- 0x3419
		"10000000",	-- 0x341a
		"10011000",	-- 0x341b
		"00000100",	-- 0x341c
		"11001100",	-- 0x341d
		"11111111",	-- 0x341e
		"01000110",	-- 0x341f
		"00000010",	-- 0x3420
		"01010010",	-- 0x3421
		"01010011",	-- 0x3422
		"01101110",	-- 0x3423
		"00101110",	-- 0x3424
		"10100111",	-- 0x3425
		"00000010",	-- 0x3426
		"01000100",	-- 0x3427
		"00000011",	-- 0x3428
		"10000110",	-- 0x3429
		"11111111",	-- 0x342a
		"11111111",	-- 0x342b
		"01101000",	-- 0x342c
		"00101110",	-- 0x342d
		"10010110",	-- 0x342e
		"11110110",	-- 0x342f
		"10001001",	-- 0x3430
		"00111101",	-- 0x3431
		"00001001",	-- 0x3432
		"01000011",	-- 0x3433
		"00000011",	-- 0x3434
		"10000110",	-- 0x3435
		"00111101",	-- 0x3436
		"00001001",	-- 0x3437
		"00000110",	-- 0x3438
		"00000110",	-- 0x3439
		"10101001",	-- 0x343a
		"00000000",	-- 0x343b
		"01000101",	-- 0x343c
		"00000010",	-- 0x343d
		"10100110",	-- 0x343e
		"00000000",	-- 0x343f
		"01111110",	-- 0x3440
		"01111110",	-- 0x3441
		"10010111",	-- 0x3442
		"00000100",	-- 0x3443
		"10101010",	-- 0x3444
		"10000000",	-- 0x3445
		"10010110",	-- 0x3446
		"00100110",	-- 0x3447
		"11100110",	-- 0x3448
		"00000000",	-- 0x3449
		"11100011",	-- 0x344a
		"00000100",	-- 0x344b
		"10011010",	-- 0x344c
		"00100110",	-- 0x344d
		"10010110",	-- 0x344e
		"00100110",	-- 0x344f
		"11100010",	-- 0x3450
		"00000100",	-- 0x3451
		"11100111",	-- 0x3452
		"00000000",	-- 0x3453
		"10010011",	-- 0x3454
		"00100111",	-- 0x3455
		"10010010",	-- 0x3456
		"00100110",	-- 0x3457
		"01111000",	-- 0x3458
		"00000111",	-- 0x3459
		"01100011",	-- 0x345a
		"00111111",	-- 0x345b
		"11001010",	-- 0x345c
		"10011100",	-- 0x345d
		"01000000",	-- 0x345e
		"00000011",	-- 0x345f
		"00111111",	-- 0x3460
		"11001010",	-- 0x3461
		"10011111",	-- 0x3462
		"11010010",	-- 0x3463
		"01000011",	-- 0x3464
		"01000110",	-- 0x3465
		"00000101",	-- 0x3466
		"00110101",	-- 0x3467
		"10010011",	-- 0x3468
		"00000010",	-- 0x3469
		"01100101",	-- 0x346a
		"01000001",	-- 0x346b
		"01100111",	-- 0x346c
		"00111101",	-- 0x346d
		"01100011",	-- 0x346e
		"11011011",	-- 0x346f
		"10100001",	-- 0x3470
		"11111010",	-- 0x3471
		"00000001",	-- 0x3472
		"10110111",	-- 0x3473
		"01011001",	-- 0x3474
		"01000110",	-- 0x3475
		"00000100",	-- 0x3476
		"01110111",	-- 0x3477
		"00100010",	-- 0x3478
		"01000000",	-- 0x3479
		"00000110",	-- 0x347a
		"11000011",	-- 0x347b
		"00000111",	-- 0x347c
		"01000110",	-- 0x347d
		"00000101",	-- 0x347e
		"01110101",	-- 0x347f
		"00100010",	-- 0x3480
		"00000011",	-- 0x3481
		"11110101",	-- 0x3482
		"00010101",	-- 0x3483
		"01010001",	-- 0x3484
		"01000110",	-- 0x3485
		"00000011",	-- 0x3486
		"00000011",	-- 0x3487
		"11110101",	-- 0x3488
		"00001011",	-- 0x3489
		"01010001",	-- 0x348a
		"01000111",	-- 0x348b
		"00000011",	-- 0x348c
		"00000011",	-- 0x348d
		"11110101",	-- 0x348e
		"00101001",	-- 0x348f
		"00110101",	-- 0x3490
		"10110000",	-- 0x3491
		"01110101",	-- 0x3492
		"00110111",	-- 0x3493
		"01000110",	-- 0x3494
		"01110010",	-- 0x3495
		"00110101",	-- 0x3496
		"10101101",	-- 0x3497
		"01101111",	-- 0x3498
		"00110101",	-- 0x3499
		"10101001",	-- 0x349a
		"01101100",	-- 0x349b
		"01111001",	-- 0x349c
		"01111010",	-- 0x349d
		"10111110",	-- 0x349e
		"01000011",	-- 0x349f
		"01100111",	-- 0x34a0
		"01111001",	-- 0x34a1
		"01111010",	-- 0x34a2
		"11000000",	-- 0x34a3
		"01000011",	-- 0x34a4
		"01100010",	-- 0x34a5
		"01011011",	-- 0x34a6
		"00110111",	-- 0x34a7
		"10100010",	-- 0x34a8
		"00000010",	-- 0x34a9
		"11000001",	-- 0x34aa
		"00000100",	-- 0x34ab
		"00010001",	-- 0x34ac
		"00010001",	-- 0x34ad
		"00010001",	-- 0x34ae
		"00010101",	-- 0x34af
		"01001000",	-- 0x34b0
		"00011110",	-- 0x34b1
		"01000101",	-- 0x34b2
		"01001011",	-- 0x34b3
		"01111001",	-- 0x34b4
		"00111001",	-- 0x34b5
		"01011001",	-- 0x34b6
		"01000101",	-- 0x34b7
		"01001111",	-- 0x34b8
		"01111001",	-- 0x34b9
		"10010000",	-- 0x34ba
		"01011001",	-- 0x34bb
		"01000100",	-- 0x34bc
		"01001010",	-- 0x34bd
		"01111001",	-- 0x34be
		"00000011",	-- 0x34bf
		"10100111",	-- 0x34c0
		"01000100",	-- 0x34c1
		"00000100",	-- 0x34c2
		"01110110",	-- 0x34c3
		"10100111",	-- 0x34c4
		"01000000",	-- 0x34c5
		"01000001",	-- 0x34c6
		"00110111",	-- 0x34c7
		"11111000",	-- 0x34c8
		"00111110",	-- 0x34c9
		"01110111",	-- 0x34ca
		"10110110",	-- 0x34cb
		"01110111",	-- 0x34cc
		"00011100",	-- 0x34cd
		"01000000",	-- 0x34ce
		"00111000",	-- 0x34cf
		"01111001",	-- 0x34d0
		"00001110",	-- 0x34d1
		"01011001",	-- 0x34d2
		"01000101",	-- 0x34d3
		"00110011",	-- 0x34d4
		"01111001",	-- 0x34d5
		"10010000",	-- 0x34d6
		"01011001",	-- 0x34d7
		"01000100",	-- 0x34d8
		"00101110",	-- 0x34d9
		"11011011",	-- 0x34da
		"10000000",	-- 0x34db
		"11001111",	-- 0x34dc
		"10000000",	-- 0x34dd
		"01000110",	-- 0x34de
		"00101000",	-- 0x34df
		"11000010",	-- 0x34e0
		"11110000",	-- 0x34e1
		"11000000",	-- 0x34e2
		"00010000",	-- 0x34e3
		"11001100",	-- 0x34e4
		"11000000",	-- 0x34e5
		"01000101",	-- 0x34e6
		"00000101",	-- 0x34e7
		"01110111",	-- 0x34e8
		"10011000",	-- 0x34e9
		"01010010",	-- 0x34ea
		"01000000",	-- 0x34eb
		"00000100",	-- 0x34ec
		"11001100",	-- 0x34ed
		"01100000",	-- 0x34ee
		"01000110",	-- 0x34ef
		"00011000",	-- 0x34f0
		"01110101",	-- 0x34f1
		"01000110",	-- 0x34f2
		"10000101",	-- 0x34f3
		"00000000",	-- 0x34f4
		"10000101",	-- 0x34f5
		"00000000",	-- 0x34f6
		"10000101",	-- 0x34f7
		"00000000",	-- 0x34f8
		"01110111",	-- 0x34f9
		"01000110",	-- 0x34fa
		"01110111",	-- 0x34fb
		"10110110",	-- 0x34fc
		"01000000",	-- 0x34fd
		"00001010",	-- 0x34fe
		"00110101",	-- 0x34ff
		"00011100",	-- 0x3500
		"00000110",	-- 0x3501
		"01110101",	-- 0x3502
		"10110110",	-- 0x3503
		"01110101",	-- 0x3504
		"10011000",	-- 0x3505
		"01110010",	-- 0x3506
		"10100111",	-- 0x3507
		"01010010",	-- 0x3508
		"01000000",	-- 0x3509
		"00011011",	-- 0x350a
		"01110101",	-- 0x350b
		"00100010",	-- 0x350c
		"01000000",	-- 0x350d
		"00000010",	-- 0x350e
		"01110111",	-- 0x350f
		"00100010",	-- 0x3510
		"01110111",	-- 0x3511
		"00000010",	-- 0x3512
		"01000000",	-- 0x3513
		"00010100",	-- 0x3514
		"00110111",	-- 0x3515
		"10100010",	-- 0x3516
		"00000010",	-- 0x3517
		"11000110",	-- 0x3518
		"00001000",	-- 0x3519
		"01110101",	-- 0x351a
		"00000010",	-- 0x351b
		"00110101",	-- 0x351c
		"10000010",	-- 0x351d
		"00000010",	-- 0x351e
		"11000110",	-- 0x351f
		"00000010",	-- 0x3520
		"00110101",	-- 0x3521
		"01100010",	-- 0x3522
		"00000010",	-- 0x3523
		"11000110",	-- 0x3524
		"00000001",	-- 0x3525
		"10110010",	-- 0x3526
		"00000001",	-- 0x3527
		"10110111",	-- 0x3528
		"01100011",	-- 0x3529
		"11011011",	-- 0x352a
		"10100010",	-- 0x352b
		"01001010",	-- 0x352c
		"00000011",	-- 0x352d
		"00000011",	-- 0x352e
		"11110110",	-- 0x352f
		"11000100",	-- 0x3530
		"11000011",	-- 0x3531
		"00001111",	-- 0x3532
		"01000110",	-- 0x3533
		"00000010",	-- 0x3534
		"01000000",	-- 0x3535
		"00000111",	-- 0x3536
		"11001101",	-- 0x3537
		"00000001",	-- 0x3538
		"01000110",	-- 0x3539
		"00000000",	-- 0x353a
		"00000011",	-- 0x353b
		"11110110",	-- 0x353c
		"11000100",	-- 0x353d
		"11111010",	-- 0x353e
		"00000001",	-- 0x353f
		"10111000",	-- 0x3540
		"01010110",	-- 0x3541
		"01000111",	-- 0x3542
		"00000011",	-- 0x3543
		"10110010",	-- 0x3544
		"00000001",	-- 0x3545
		"10111000",	-- 0x3546
		"11011010",	-- 0x3547
		"01011001",	-- 0x3548
		"11001100",	-- 0x3549
		"10010000",	-- 0x354a
		"01000100",	-- 0x354b
		"00011101",	-- 0x354c
		"11001100",	-- 0x354d
		"00010000",	-- 0x354e
		"01000101",	-- 0x354f
		"00100010",	-- 0x3550
		"00110101",	-- 0x3551
		"01010110",	-- 0x3552
		"00011111",	-- 0x3553
		"11111010",	-- 0x3554
		"00000010",	-- 0x3555
		"00111010",	-- 0x3556
		"11001100",	-- 0x3557
		"00000100",	-- 0x3558
		"01000101",	-- 0x3559
		"00011000",	-- 0x355a
		"01111001",	-- 0x355b
		"11010010",	-- 0x355c
		"01010111",	-- 0x355d
		"01000101",	-- 0x355e
		"00010011",	-- 0x355f
		"01110111",	-- 0x3560
		"11111000",	-- 0x3561
		"00110111",	-- 0x3562
		"10110110",	-- 0x3563
		"00010111",	-- 0x3564
		"11111010",	-- 0x3565
		"00000001",	-- 0x3566
		"10111001",	-- 0x3567
		"01000000",	-- 0x3568
		"00001101",	-- 0x3569
		"00110111",	-- 0x356a
		"11111000",	-- 0x356b
		"00000110",	-- 0x356c
		"11111010",	-- 0x356d
		"00000001",	-- 0x356e
		"10110011",	-- 0x356f
		"10110010",	-- 0x3570
		"00000001",	-- 0x3571
		"10110101",	-- 0x3572
		"01110101",	-- 0x3573
		"11111000",	-- 0x3574
		"11001010",	-- 0x3575
		"00011010",	-- 0x3576
		"01110010",	-- 0x3577
		"11100011",	-- 0x3578
		"00000011",	-- 0x3579
		"11110110",	-- 0x357a
		"00000000",	-- 0x357b
		"11111010",	-- 0x357c
		"00000001",	-- 0x357d
		"10110111",	-- 0x357e
		"11000010",	-- 0x357f
		"00000011",	-- 0x3580
		"01000111",	-- 0x3581
		"00111010",	-- 0x3582
		"10001111",	-- 0x3583
		"11000011",	-- 0x3584
		"10010100",	-- 0x3585
		"00001101",	-- 0x3586
		"11101010",	-- 0x3587
		"10000000",	-- 0x3588
		"11111011",	-- 0x3589
		"00000001",	-- 0x358a
		"10111000",	-- 0x358b
		"11001101",	-- 0x358c
		"00000100",	-- 0x358d
		"01000010",	-- 0x358e
		"00001101",	-- 0x358f
		"00010010",	-- 0x3590
		"11001101",	-- 0x3591
		"00000001",	-- 0x3592
		"01000010",	-- 0x3593
		"00001000",	-- 0x3594
		"01101101",	-- 0x3595
		"11111011",	-- 0x3596
		"00000010",	-- 0x3597
		"00010110",	-- 0x3598
		"01111101",	-- 0x3599
		"01000110",	-- 0x359a
		"00000001",	-- 0x359b
		"00010010",	-- 0x359c
		"11110000",	-- 0x359d
		"00000001",	-- 0x359e
		"10110011",	-- 0x359f
		"01000100",	-- 0x35a0
		"00000010",	-- 0x35a1
		"11001010",	-- 0x35a2
		"11111111",	-- 0x35a3
		"10110010",	-- 0x35a4
		"00000001",	-- 0x35a5
		"10110011",	-- 0x35a6
		"11001101",	-- 0x35a7
		"00000100",	-- 0x35a8
		"01000101",	-- 0x35a9
		"00001110",	-- 0x35aa
		"11110100",	-- 0x35ab
		"00000001",	-- 0x35ac
		"10111010",	-- 0x35ad
		"01000011",	-- 0x35ae
		"00001001",	-- 0x35af
		"00010000",	-- 0x35b0
		"00010000",	-- 0x35b1
		"01010110",	-- 0x35b2
		"11110000",	-- 0x35b3
		"00000001",	-- 0x35b4
		"10111010",	-- 0x35b5
		"10110010",	-- 0x35b6
		"00000001",	-- 0x35b7
		"10111010",	-- 0x35b8
		"01010010",	-- 0x35b9
		"10110010",	-- 0x35ba
		"00000001",	-- 0x35bb
		"10111000",	-- 0x35bc
		"11111010",	-- 0x35bd
		"00000001",	-- 0x35be
		"10111001",	-- 0x35bf
		"01011011",	-- 0x35c0
		"11110100",	-- 0x35c1
		"00000001",	-- 0x35c2
		"10111011",	-- 0x35c3
		"01000100",	-- 0x35c4
		"00001000",	-- 0x35c5
		"11110000",	-- 0x35c6
		"00000001",	-- 0x35c7
		"10110011",	-- 0x35c8
		"01000101",	-- 0x35c9
		"00001000",	-- 0x35ca
		"01010010",	-- 0x35cb
		"01000000",	-- 0x35cc
		"00000101",	-- 0x35cd
		"11110000",	-- 0x35ce
		"00000001",	-- 0x35cf
		"10110011",	-- 0x35d0
		"01000101",	-- 0x35d1
		"00000011",	-- 0x35d2
		"00001011",	-- 0x35d3
		"01000011",	-- 0x35d4
		"00000001",	-- 0x35d5
		"01011010",	-- 0x35d6
		"11111011",	-- 0x35d7
		"00000001",	-- 0x35d8
		"01010111",	-- 0x35d9
		"00010011",	-- 0x35da
		"01000101",	-- 0x35db
		"00010111",	-- 0x35dc
		"11110101",	-- 0x35dd
		"00000010",	-- 0x35de
		"00111010",	-- 0x35df
		"01000100",	-- 0x35e0
		"00010010",	-- 0x35e1
		"11110001",	-- 0x35e2
		"00000001",	-- 0x35e3
		"10111001",	-- 0x35e4
		"01000101",	-- 0x35e5
		"00000001",	-- 0x35e6
		"01010011",	-- 0x35e7
		"00001011",	-- 0x35e8
		"01000011",	-- 0x35e9
		"00001001",	-- 0x35ea
		"01011010",	-- 0x35eb
		"11001100",	-- 0x35ec
		"00011010",	-- 0x35ed
		"01000100",	-- 0x35ee
		"00000010",	-- 0x35ef
		"11001010",	-- 0x35f0
		"00011010",	-- 0x35f1
		"01000000",	-- 0x35f2
		"00001100",	-- 0x35f3
		"11111011",	-- 0x35f4
		"00000001",	-- 0x35f5
		"01101000",	-- 0x35f6
		"01000110",	-- 0x35f7
		"00000111",	-- 0x35f8
		"11111100",	-- 0x35f9
		"00000001",	-- 0x35fa
		"10111010",	-- 0x35fb
		"01000010",	-- 0x35fc
		"00000111",	-- 0x35fd
		"01011011",	-- 0x35fe
		"10001100",	-- 0x35ff
		"11001011",	-- 0x3600
		"00011010",	-- 0x3601
		"10110011",	-- 0x3602
		"00000001",	-- 0x3603
		"10111010",	-- 0x3604
		"10110010",	-- 0x3605
		"00000001",	-- 0x3606
		"10110011",	-- 0x3607
		"11111010",	-- 0x3608
		"00000001",	-- 0x3609
		"10111001",	-- 0x360a
		"10110010",	-- 0x360b
		"00000001",	-- 0x360c
		"10111011",	-- 0x360d
		"01010010",	-- 0x360e
		"00110101",	-- 0x360f
		"01010110",	-- 0x3610
		"00101111",	-- 0x3611
		"11111010",	-- 0x3612
		"00000001",	-- 0x3613
		"10110011",	-- 0x3614
		"01111001",	-- 0x3615
		"11010010",	-- 0x3616
		"01010111",	-- 0x3617
		"01000100",	-- 0x3618
		"00000100",	-- 0x3619
		"11000000",	-- 0x361a
		"00000000",	-- 0x361b
		"01000000",	-- 0x361c
		"00010011",	-- 0x361d
		"11001011",	-- 0x361e
		"10010000",	-- 0x361f
		"11001101",	-- 0x3620
		"10010001",	-- 0x3621
		"01000100",	-- 0x3622
		"00001101",	-- 0x3623
		"01111001",	-- 0x3624
		"10010000",	-- 0x3625
		"01011001",	-- 0x3626
		"01000101",	-- 0x3627
		"00001000",	-- 0x3628
		"11111010",	-- 0x3629
		"00000001",	-- 0x362a
		"10110101",	-- 0x362b
		"11110100",	-- 0x362c
		"00000011",	-- 0x362d
		"00000110",	-- 0x362e
		"01000000",	-- 0x362f
		"00000011",	-- 0x3630
		"11110100",	-- 0x3631
		"00000001",	-- 0x3632
		"10111001",	-- 0x3633
		"01000100",	-- 0x3634
		"00001000",	-- 0x3635
		"11110000",	-- 0x3636
		"00000010",	-- 0x3637
		"00111010",	-- 0x3638
		"01000101",	-- 0x3639
		"00000110",	-- 0x363a
		"01010010",	-- 0x363b
		"01000000",	-- 0x363c
		"00000011",	-- 0x363d
		"11111010",	-- 0x363e
		"00000010",	-- 0x363f
		"00111010",	-- 0x3640
		"10110010",	-- 0x3641
		"00000010",	-- 0x3642
		"00010110",	-- 0x3643
		"01111001",	-- 0x3644
		"01000000",	-- 0x3645
		"11001011",	-- 0x3646
		"01000100",	-- 0x3647
		"00000011",	-- 0x3648
		"00000011",	-- 0x3649
		"11110110",	-- 0x364a
		"11000100",	-- 0x364b
		"01110010",	-- 0x364c
		"11001011",	-- 0x364d
		"11111010",	-- 0x364e
		"00000001",	-- 0x364f
		"10110011",	-- 0x3650
		"11000100",	-- 0x3651
		"00000010",	-- 0x3652
		"01000100",	-- 0x3653
		"00000001",	-- 0x3654
		"01010010",	-- 0x3655
		"11111011",	-- 0x3656
		"00000010",	-- 0x3657
		"00010110",	-- 0x3658
		"01000110",	-- 0x3659
		"00000110",	-- 0x365a
		"11001100",	-- 0x365b
		"00011010",	-- 0x365c
		"01000100",	-- 0x365d
		"00000010",	-- 0x365e
		"11001010",	-- 0x365f
		"00011010",	-- 0x3660
		"10110010",	-- 0x3661
		"00000001",	-- 0x3662
		"10110011",	-- 0x3663
		"11111011",	-- 0x3664
		"00000001",	-- 0x3665
		"10111001",	-- 0x3666
		"01000111",	-- 0x3667
		"00111010",	-- 0x3668
		"11011010",	-- 0x3669
		"01011001",	-- 0x366a
		"11001100",	-- 0x366b
		"00011000",	-- 0x366c
		"01000101",	-- 0x366d
		"00110100",	-- 0x366e
		"11001100",	-- 0x366f
		"10001100",	-- 0x3670
		"01000100",	-- 0x3671
		"00110000",	-- 0x3672
		"11111010",	-- 0x3673
		"00000001",	-- 0x3674
		"10111010",	-- 0x3675
		"11000100",	-- 0x3676
		"00010001",	-- 0x3677
		"01000100",	-- 0x3678
		"00010010",	-- 0x3679
		"11111010",	-- 0x367a
		"00000001",	-- 0x367b
		"10111100",	-- 0x367c
		"10001111",	-- 0x367d
		"11000011",	-- 0x367e
		"10011000",	-- 0x367f
		"00001101",	-- 0x3680
		"11101010",	-- 0x3681
		"10000000",	-- 0x3682
		"00001000",	-- 0x3683
		"11001100",	-- 0x3684
		"10101011",	-- 0x3685
		"01000011",	-- 0x3686
		"00000010",	-- 0x3687
		"11001010",	-- 0x3688
		"10101011",	-- 0x3689
		"01000000",	-- 0x368a
		"00001110",	-- 0x368b
		"11000100",	-- 0x368c
		"00010001",	-- 0x368d
		"01000011",	-- 0x368e
		"00010011",	-- 0x368f
		"00000010",	-- 0x3690
		"00001001",	-- 0x3691
		"01000101",	-- 0x3692
		"00000100",	-- 0x3693
		"11001100",	-- 0x3694
		"00011010",	-- 0x3695
		"01000100",	-- 0x3696
		"00000010",	-- 0x3697
		"11001010",	-- 0x3698
		"00011010",	-- 0x3699
		"10001111",	-- 0x369a
		"00000011",	-- 0x369b
		"00000100",	-- 0x369c
		"11111011",	-- 0x369d
		"00000001",	-- 0x369e
		"10111100",	-- 0x369f
		"00001111",	-- 0x36a0
		"10100010",	-- 0x36a1
		"10000000",	-- 0x36a2
		"10001110",	-- 0x36a3
		"11000011",	-- 0x36a4
		"10011011",	-- 0x36a5
		"11111011",	-- 0x36a6
		"00000001",	-- 0x36a7
		"10111100",	-- 0x36a8
		"00010011",	-- 0x36a9
		"00001110",	-- 0x36aa
		"11011010",	-- 0x36ab
		"01011011",	-- 0x36ac
		"01010011",	-- 0x36ad
		"11101100",	-- 0x36ae
		"00000000",	-- 0x36af
		"01000101",	-- 0x36b0
		"00000110",	-- 0x36b1
		"01010111",	-- 0x36b2
		"11101100",	-- 0x36b3
		"00000001",	-- 0x36b4
		"01000101",	-- 0x36b5
		"00000001",	-- 0x36b6
		"01010111",	-- 0x36b7
		"10110011",	-- 0x36b8
		"00000001",	-- 0x36b9
		"10111100",	-- 0x36ba
		"10001111",	-- 0x36bb
		"00000011",	-- 0x36bc
		"00000100",	-- 0x36bd
		"00001111",	-- 0x36be
		"11101010",	-- 0x36bf
		"10000000",	-- 0x36c0
		"10110010",	-- 0x36c1
		"00000001",	-- 0x36c2
		"10111001",	-- 0x36c3
		"01100011",	-- 0x36c4
		"00110111",	-- 0x36c5
		"10110110",	-- 0x36c6
		"00001011",	-- 0x36c7
		"00000101",	-- 0x36c8
		"10000110",	-- 0x36c9
		"10011010",	-- 0x36ca
		"10011010",	-- 0x36cb
		"10111010",	-- 0x36cc
		"00000011",	-- 0x36cd
		"00000100",	-- 0x36ce
		"10110010",	-- 0x36cf
		"00000011",	-- 0x36d0
		"00000110",	-- 0x36d1
		"00000111",	-- 0x36d2
		"01111001",	-- 0x36d3
		"11010010",	-- 0x36d4
		"01010111",	-- 0x36d5
		"01000101",	-- 0x36d6
		"00001101",	-- 0x36d7
		"00110101",	-- 0x36d8
		"10110110",	-- 0x36d9
		"00001010",	-- 0x36da
		"11011010",	-- 0x36db
		"01011100",	-- 0x36dc
		"11001100",	-- 0x36dd
		"10010110",	-- 0x36de
		"01000100",	-- 0x36df
		"00000110",	-- 0x36e0
		"11001100",	-- 0x36e1
		"01101010",	-- 0x36e2
		"01000011",	-- 0x36e3
		"00000010",	-- 0x36e4
		"01110010",	-- 0x36e5
		"11001100",	-- 0x36e6
		"01111001",	-- 0x36e7
		"00000110",	-- 0x36e8
		"11001100",	-- 0x36e9
		"01000101",	-- 0x36ea
		"00000011",	-- 0x36eb
		"01110111",	-- 0x36ec
		"01000010",	-- 0x36ed
		"10001100",	-- 0x36ee
		"01110101",	-- 0x36ef
		"01000010",	-- 0x36f0
		"01100011",	-- 0x36f1
		"01101110",	-- 0x36f2
		"01101111",	-- 0x36f3
		"01110101",	-- 0x36f4
		"00001100",	-- 0x36f5
		"00110111",	-- 0x36f6
		"00000101",	-- 0x36f7
		"01111001",	-- 0x36f8
		"01110101",	-- 0x36f9
		"00010101",	-- 0x36fa
		"00110111",	-- 0x36fb
		"10110101",	-- 0x36fc
		"00000111",	-- 0x36fd
		"01110101",	-- 0x36fe
		"10110101",	-- 0x36ff
		"00000001",	-- 0x3700
		"11110010",	-- 0x3701
		"01001011",	-- 0x3702
		"01000000",	-- 0x3703
		"00001011",	-- 0x3704
		"10010110",	-- 0x3705
		"00001000",	-- 0x3706
		"10000111",	-- 0x3707
		"00111111",	-- 0x3708
		"01111010",	-- 0x3709
		"10011010",	-- 0x370a
		"00001000",	-- 0x370b
		"01110101",	-- 0x370c
		"00000110",	-- 0x370d
		"01110111",	-- 0x370e
		"00110101",	-- 0x370f
		"01110001",	-- 0x3710
		"01110101",	-- 0x3711
		"01000110",	-- 0x3712
		"01011100",	-- 0x3713
		"00000001",	-- 0x3714
		"11011101",	-- 0x3715
		"01010011",	-- 0x3716
		"00110101",	-- 0x3717
		"10001101",	-- 0x3718
		"00111000",	-- 0x3719
		"10110110",	-- 0x371a
		"00000001",	-- 0x371b
		"10001010",	-- 0x371c
		"01010110",	-- 0x371d
		"01000110",	-- 0x371e
		"00000001",	-- 0x371f
		"01010000",	-- 0x3720
		"11001100",	-- 0x3721
		"00000101",	-- 0x3722
		"01000101",	-- 0x3723
		"00000010",	-- 0x3724
		"01110111",	-- 0x3725
		"10010011",	-- 0x3726
		"01111001",	-- 0x3727
		"00111111",	-- 0x3728
		"11000010",	-- 0x3729
		"01000101",	-- 0x372a
		"00101110",	-- 0x372b
		"01111001",	-- 0x372c
		"00111100",	-- 0x372d
		"01011001",	-- 0x372e
		"01000101",	-- 0x372f
		"00001000",	-- 0x3730
		"01111001",	-- 0x3731
		"01110011",	-- 0x3732
		"01010110",	-- 0x3733
		"01000101",	-- 0x3734
		"00100100",	-- 0x3735
		"00110101",	-- 0x3736
		"00011001",	-- 0x3737
		"00100001",	-- 0x3738
		"11001101",	-- 0x3739
		"00000001",	-- 0x373a
		"01000010",	-- 0x373b
		"00000010",	-- 0x373c
		"01110010",	-- 0x373d
		"11000001",	-- 0x373e
		"01010111",	-- 0x373f
		"01000110",	-- 0x3740
		"00000001",	-- 0x3741
		"01010001",	-- 0x3742
		"11001101",	-- 0x3743
		"00001001",	-- 0x3744
		"01000101",	-- 0x3745
		"00010101",	-- 0x3746
		"01111001",	-- 0x3747
		"00111111",	-- 0x3748
		"11000001",	-- 0x3749
		"01000101",	-- 0x374a
		"00010000",	-- 0x374b
		"01110111",	-- 0x374c
		"01011011",	-- 0x374d
		"01110111",	-- 0x374e
		"10011101",	-- 0x374f
		"01000000",	-- 0x3750
		"00001010",	-- 0x3751
		"01110101",	-- 0x3752
		"10001101",	-- 0x3753
		"01110101",	-- 0x3754
		"10010011",	-- 0x3755
		"01110101",	-- 0x3756
		"01011011",	-- 0x3757
		"11001010",	-- 0x3758
		"00000001",	-- 0x3759
		"11001011",	-- 0x375a
		"00000001",	-- 0x375b
		"10111010",	-- 0x375c
		"00000001",	-- 0x375d
		"10001010",	-- 0x375e
		"01000000",	-- 0x375f
		"00001111",	-- 0x3760
		"00110101",	-- 0x3761
		"10011101",	-- 0x3762
		"00000010",	-- 0x3763
		"01110010",	-- 0x3764
		"11100111",	-- 0x3765
		"11000010",	-- 0x3766
		"11111011",	-- 0x3767
		"01111001",	-- 0x3768
		"00101110",	-- 0x3769
		"11100111",	-- 0x376a
		"01000011",	-- 0x376b
		"00000010",	-- 0x376c
		"11000110",	-- 0x376d
		"00000100",	-- 0x376e
		"01100011",	-- 0x376f
		"01000000",	-- 0x3770
		"00100101",	-- 0x3771
		"10010110",	-- 0x3772
		"00001000",	-- 0x3773
		"10111010",	-- 0x3774
		"00000001",	-- 0x3775
		"01110000",	-- 0x3776
		"00110101",	-- 0x3777
		"10110000",	-- 0x3778
		"00000110",	-- 0x3779
		"00110101",	-- 0x377a
		"00011001",	-- 0x377b
		"00000011",	-- 0x377c
		"01110101",	-- 0x377d
		"01010101",	-- 0x377e
		"10001100",	-- 0x377f
		"01110111",	-- 0x3780
		"01010101",	-- 0x3781
		"00110111",	-- 0x3782
		"01110101",	-- 0x3783
		"00000100",	-- 0x3784
		"01110101",	-- 0x3785
		"01110101",	-- 0x3786
		"01110111",	-- 0x3787
		"10010101",	-- 0x3788
		"00110101",	-- 0x3789
		"00110101",	-- 0x378a
		"00001011",	-- 0x378b
		"00110101",	-- 0x378c
		"01010101",	-- 0x378d
		"00001000",	-- 0x378e
		"10010110",	-- 0x378f
		"11110110",	-- 0x3790
		"10110111",	-- 0x3791
		"00000001",	-- 0x3792
		"01110000",	-- 0x3793
		"00000001",	-- 0x3794
		"11110010",	-- 0x3795
		"00001001",	-- 0x3796
		"01111111",	-- 0x3797
		"01111110",	-- 0x3798
		"01110011",	-- 0x3799
		"01110101",	-- 0x379a
		"10001100",	-- 0x379b
		"01101110",	-- 0x379c
		"01101111",	-- 0x379d
		"11011010",	-- 0x379e
		"11111110",	-- 0x379f
		"01011011",	-- 0x37a0
		"11000011",	-- 0x37a1
		"00000011",	-- 0x37a2
		"01000111",	-- 0x37a3
		"00000101",	-- 0x37a4
		"11000000",	-- 0x37a5
		"10000000",	-- 0x37a6
		"01000100",	-- 0x37a7
		"00001011",	-- 0x37a8
		"01010010",	-- 0x37a9
		"11001011",	-- 0x37aa
		"00000000",	-- 0x37ab
		"10010011",	-- 0x37ac
		"11111101",	-- 0x37ad
		"01110111",	-- 0x37ae
		"00101011",	-- 0x37af
		"01100111",	-- 0x37b0
		"00010111",	-- 0x37b1
		"10010011",	-- 0x37b2
		"00000110",	-- 0x37b3
		"10010010",	-- 0x37b4
		"11111110",	-- 0x37b5
		"00000001",	-- 0x37b6
		"11010011",	-- 0x37b7
		"10001001",	-- 0x37b8
		"11011010",	-- 0x37b9
		"00000100",	-- 0x37ba
		"00010000",	-- 0x37bb
		"00010000",	-- 0x37bc
		"00010000",	-- 0x37bd
		"01000100",	-- 0x37be
		"00000000",	-- 0x37bf
		"01110101",	-- 0x37c0
		"01010010",	-- 0x37c1
		"01110111",	-- 0x37c2
		"00101101",	-- 0x37c3
		"01111111",	-- 0x37c4
		"01111110",	-- 0x37c5
		"01110011",	-- 0x37c6
		"10000110",	-- 0x37c7
		"10101101",	-- 0x37c8
		"00011001",	-- 0x37c9
		"00000001",	-- 0x37ca
		"11000100",	-- 0x37cb
		"10111001",	-- 0x37cc
		"00000001",	-- 0x37cd
		"11111011",	-- 0x37ce
		"00011101",	-- 0x37cf
		"11011011",	-- 0x37d0
		"10101011",	-- 0x37d1
		"01110001",	-- 0x37d2
		"01100110",	-- 0x37d3
		"01000111",	-- 0x37d4
		"01000111",	-- 0x37d5
		"11111010",	-- 0x37d6
		"00000010",	-- 0x37d7
		"01000010",	-- 0x37d8
		"11001110",	-- 0x37d9
		"00000100",	-- 0x37da
		"01000111",	-- 0x37db
		"00000111",	-- 0x37dc
		"00110101",	-- 0x37dd
		"01110111",	-- 0x37de
		"00011101",	-- 0x37df
		"01110111",	-- 0x37e0
		"01110111",	-- 0x37e1
		"01000000",	-- 0x37e2
		"00000101",	-- 0x37e3
		"00110111",	-- 0x37e4
		"01110111",	-- 0x37e5
		"00010110",	-- 0x37e6
		"01110101",	-- 0x37e7
		"01110111",	-- 0x37e8
		"01110010",	-- 0x37e9
		"10101100",	-- 0x37ea
		"11000001",	-- 0x37eb
		"00010000",	-- 0x37ec
		"11001101",	-- 0x37ed
		"00100000",	-- 0x37ee
		"01000101",	-- 0x37ef
		"00101010",	-- 0x37f0
		"11001011",	-- 0x37f1
		"00100000",	-- 0x37f2
		"11011010",	-- 0x37f3
		"01101101",	-- 0x37f4
		"11000010",	-- 0x37f5
		"11111110",	-- 0x37f6
		"10010010",	-- 0x37f7
		"01101101",	-- 0x37f8
		"01110101",	-- 0x37f9
		"11110110",	-- 0x37fa
		"01000000",	-- 0x37fb
		"00011110",	-- 0x37fc
		"01110110",	-- 0x37fd
		"10101100",	-- 0x37fe
		"01111001",	-- 0x37ff
		"00010110",	-- 0x3800
		"10101100",	-- 0x3801
		"01000101",	-- 0x3802
		"00010111",	-- 0x3803
		"01110101",	-- 0x3804
		"01110111",	-- 0x3805
		"01110101",	-- 0x3806
		"01100110",	-- 0x3807
		"01110010",	-- 0x3808
		"10101100",	-- 0x3809
		"11000011",	-- 0x380a
		"00001111",	-- 0x380b
		"01010111",	-- 0x380c
		"11001101",	-- 0x380d
		"00000011",	-- 0x380e
		"01000101",	-- 0x380f
		"00001010",	-- 0x3810
		"11001011",	-- 0x3811
		"00000011",	-- 0x3812
		"11011010",	-- 0x3813
		"01101101",	-- 0x3814
		"11000110",	-- 0x3815
		"00000001",	-- 0x3816
		"10010010",	-- 0x3817
		"01101101",	-- 0x3818
		"01110111",	-- 0x3819
		"11110110",	-- 0x381a
		"10010011",	-- 0x381b
		"10101011",	-- 0x381c
		"00000001",	-- 0x381d
		"11111000",	-- 0x381e
		"01111100",	-- 0x381f
		"00000001",	-- 0x3820
		"11110000",	-- 0x3821
		"00110011",	-- 0x3822
		"00000001",	-- 0x3823
		"11101011",	-- 0x3824
		"11110011",	-- 0x3825
		"01110110",	-- 0x3826
		"11000110",	-- 0x3827
		"11001010",	-- 0x3828
		"00000001",	-- 0x3829
		"11011110",	-- 0x382a
		"11000110",	-- 0x382b
		"01000111",	-- 0x382c
		"00000011",	-- 0x382d
		"00000001",	-- 0x382e
		"11100111",	-- 0x382f
		"10011110",	-- 0x3830
		"00000001",	-- 0x3831
		"11100111",	-- 0x3832
		"10110001",	-- 0x3833
		"01111001",	-- 0x3834
		"01010110",	-- 0x3835
		"10110010",	-- 0x3836
		"01000101",	-- 0x3837
		"00010100",	-- 0x3838
		"01110010",	-- 0x3839
		"10110010",	-- 0x383a
		"00000001",	-- 0x383b
		"11001100",	-- 0x383c
		"10110111",	-- 0x383d
		"00000001",	-- 0x383e
		"11111001",	-- 0x383f
		"11101101",	-- 0x3840
		"10010110",	-- 0x3841
		"01011001",	-- 0x3842
		"00000100",	-- 0x3843
		"00000100",	-- 0x3844
		"10010101",	-- 0x3845
		"01011101",	-- 0x3846
		"01000100",	-- 0x3847
		"00000010",	-- 0x3848
		"11001011",	-- 0x3849
		"11111111",	-- 0x384a
		"10010011",	-- 0x384b
		"11111011",	-- 0x384c
		"00110111",	-- 0x384d
		"00110010",	-- 0x384e
		"00101001",	-- 0x384f
		"11011010",	-- 0x3850
		"00000100",	-- 0x3851
		"00010000",	-- 0x3852
		"00010000",	-- 0x3853
		"00010000",	-- 0x3854
		"01000101",	-- 0x3855
		"00011001",	-- 0x3856
		"00010000",	-- 0x3857
		"01000101",	-- 0x3858
		"00010000",	-- 0x3859
		"00010000",	-- 0x385a
		"01000101",	-- 0x385b
		"00001001",	-- 0x385c
		"00010000",	-- 0x385d
		"01000101",	-- 0x385e
		"00000010",	-- 0x385f
		"01000000",	-- 0x3860
		"00010111",	-- 0x3861
		"01110101",	-- 0x3862
		"11110001",	-- 0x3863
		"01000000",	-- 0x3864
		"00010011",	-- 0x3865
		"01110101",	-- 0x3866
		"11010001",	-- 0x3867
		"01000000",	-- 0x3868
		"00001111",	-- 0x3869
		"01110101",	-- 0x386a
		"10110001",	-- 0x386b
		"01110101",	-- 0x386c
		"10010001",	-- 0x386d
		"01000000",	-- 0x386e
		"00001001",	-- 0x386f
		"10000110",	-- 0x3870
		"11000111",	-- 0x3871
		"00000110",	-- 0x3872
		"00000001",	-- 0x3873
		"11000100",	-- 0x3874
		"10111001",	-- 0x3875
		"00000001",	-- 0x3876
		"11111001",	-- 0x3877
		"00100010",	-- 0x3878
		"01110111",	-- 0x3879
		"11110010",	-- 0x387a
		"01100011",	-- 0x387b
		"01111001",	-- 0x387c
		"00000100",	-- 0x387d
		"11000101",	-- 0x387e
		"01000011",	-- 0x387f
		"00001100",	-- 0x3880
		"11111010",	-- 0x3881
		"00000001",	-- 0x3882
		"11011101",	-- 0x3883
		"11000010",	-- 0x3884
		"10111111",	-- 0x3885
		"10110010",	-- 0x3886
		"00000001",	-- 0x3887
		"11011101",	-- 0x3888
		"10010010",	-- 0x3889
		"00010010",	-- 0x388a
		"01000000",	-- 0x388b
		"00001010",	-- 0x388c
		"11011010",	-- 0x388d
		"00000011",	-- 0x388e
		"11001110",	-- 0x388f
		"01000000",	-- 0x3890
		"01000111",	-- 0x3891
		"00011000",	-- 0x3892
		"11001110",	-- 0x3893
		"00001000",	-- 0x3894
		"01000110",	-- 0x3895
		"00000010",	-- 0x3896
		"01110010",	-- 0x3897
		"11000101",	-- 0x3898
		"11111010",	-- 0x3899
		"00000001",	-- 0x389a
		"11011101",	-- 0x389b
		"11000110",	-- 0x389c
		"01000000",	-- 0x389d
		"10110010",	-- 0x389e
		"00000001",	-- 0x389f
		"11011101",	-- 0x38a0
		"10010010",	-- 0x38a1
		"00010010",	-- 0x38a2
		"10000110",	-- 0x38a3
		"10010010",	-- 0x38a4
		"00000000",	-- 0x38a5
		"10011010",	-- 0x38a6
		"00011010",	-- 0x38a7
		"00110011",	-- 0x38a8
		"10110111",	-- 0x38a9
		"00000011",	-- 0x38aa
		"01111001",	-- 0x38ab
		"00100100",	-- 0x38ac
		"01110110",	-- 0x38ad
		"01000101",	-- 0x38ae
		"00010100",	-- 0x38af
		"01110101",	-- 0x38b0
		"01001111",	-- 0x38b1
		"11111010",	-- 0x38b2
		"00000001",	-- 0x38b3
		"11011101",	-- 0x38b4
		"11000010",	-- 0x38b5
		"01111111",	-- 0x38b6
		"10110010",	-- 0x38b7
		"00000001",	-- 0x38b8
		"11011101",	-- 0x38b9
		"10010010",	-- 0x38ba
		"00010010",	-- 0x38bb
		"11011010",	-- 0x38bc
		"00000011",	-- 0x38bd
		"11000110",	-- 0x38be
		"10000000",	-- 0x38bf
		"10010010",	-- 0x38c0
		"00000011",	-- 0x38c1
		"01000000",	-- 0x38c2
		"00101001",	-- 0x38c3
		"01110111",	-- 0x38c4
		"01001111",	-- 0x38c5
		"01111001",	-- 0x38c6
		"00000100",	-- 0x38c7
		"11000100",	-- 0x38c8
		"01000011",	-- 0x38c9
		"00101000",	-- 0x38ca
		"11111010",	-- 0x38cb
		"00000001",	-- 0x38cc
		"11011101",	-- 0x38cd
		"11000010",	-- 0x38ce
		"01111111",	-- 0x38cf
		"10010010",	-- 0x38d0
		"00010010",	-- 0x38d1
		"11000110",	-- 0x38d2
		"10000000",	-- 0x38d3
		"10110010",	-- 0x38d4
		"00000001",	-- 0x38d5
		"11011101",	-- 0x38d6
		"10010010",	-- 0x38d7
		"00010010",	-- 0x38d8
		"10000110",	-- 0x38d9
		"10000001",	-- 0x38da
		"11011110",	-- 0x38db
		"10011010",	-- 0x38dc
		"00011000",	-- 0x38dd
		"00110011",	-- 0x38de
		"01001111",	-- 0x38df
		"00000011",	-- 0x38e0
		"11011011",	-- 0x38e1
		"01110111",	-- 0x38e2
		"01010111",	-- 0x38e3
		"01000110",	-- 0x38e4
		"00000001",	-- 0x38e5
		"01010001",	-- 0x38e6
		"10010011",	-- 0x38e7
		"01110111",	-- 0x38e8
		"11001101",	-- 0x38e9
		"00000011",	-- 0x38ea
		"01000101",	-- 0x38eb
		"00000100",	-- 0x38ec
		"01110111",	-- 0x38ed
		"11110110",	-- 0x38ee
		"01110101",	-- 0x38ef
		"01001011",	-- 0x38f0
		"01110010",	-- 0x38f1
		"11000100",	-- 0x38f2
		"01100011",	-- 0x38f3
		"01101110",	-- 0x38f4
		"01101111",	-- 0x38f5
		"01110101",	-- 0x38f6
		"01001101",	-- 0x38f7
		"11011011",	-- 0x38f8
		"01110110",	-- 0x38f9
		"11011010",	-- 0x38fa
		"00000011",	-- 0x38fb
		"11001110",	-- 0x38fc
		"00110000",	-- 0x38fd
		"01000110",	-- 0x38fe
		"00001101",	-- 0x38ff
		"00110101",	-- 0x3900
		"01001010",	-- 0x3901
		"00001010",	-- 0x3902
		"00000001",	-- 0x3903
		"11111001",	-- 0x3904
		"10011011",	-- 0x3905
		"01110010",	-- 0x3906
		"11000100",	-- 0x3907
		"01110010",	-- 0x3908
		"01110111",	-- 0x3909
		"01010011",	-- 0x390a
		"01000000",	-- 0x390b
		"00000100",	-- 0x390c
		"01010111",	-- 0x390d
		"01000110",	-- 0x390e
		"00000001",	-- 0x390f
		"01010001",	-- 0x3910
		"10010011",	-- 0x3911
		"01110110",	-- 0x3912
		"10000110",	-- 0x3913
		"10000001",	-- 0x3914
		"11011110",	-- 0x3915
		"10011010",	-- 0x3916
		"00011000",	-- 0x3917
		"00110011",	-- 0x3918
		"01001111",	-- 0x3919
		"00000011",	-- 0x391a
		"11011011",	-- 0x391b
		"00101010",	-- 0x391c
		"11011011",	-- 0x391d
		"00011100",	-- 0x391e
		"01111111",	-- 0x391f
		"01111110",	-- 0x3920
		"01110011",	-- 0x3921
		"11011010",	-- 0x3922
		"10011000",	-- 0x3923
		"00110101",	-- 0x3924
		"00010010",	-- 0x3925
		"00000010",	-- 0x3926
		"11001010",	-- 0x3927
		"01010000",	-- 0x3928
		"10110010",	-- 0x3929
		"00000010",	-- 0x392a
		"00001101",	-- 0x392b
		"11011010",	-- 0x392c
		"10010110",	-- 0x392d
		"00110101",	-- 0x392e
		"00010010",	-- 0x392f
		"00000010",	-- 0x3930
		"11001010",	-- 0x3931
		"00000000",	-- 0x3932
		"10110010",	-- 0x3933
		"00000010",	-- 0x3934
		"00010000",	-- 0x3935
		"11011010",	-- 0x3936
		"11010000",	-- 0x3937
		"10110010",	-- 0x3938
		"00000010",	-- 0x3939
		"00001110",	-- 0x393a
		"11011010",	-- 0x393b
		"11101010",	-- 0x393c
		"10110010",	-- 0x393d
		"00000010",	-- 0x393e
		"00001111",	-- 0x393f
		"11011010",	-- 0x3940
		"01100000",	-- 0x3941
		"10110010",	-- 0x3942
		"00000010",	-- 0x3943
		"00010001",	-- 0x3944
		"10110110",	-- 0x3945
		"00000001",	-- 0x3946
		"00001010",	-- 0x3947
		"10111010",	-- 0x3948
		"00000010",	-- 0x3949
		"00000110",	-- 0x394a
		"10110110",	-- 0x394b
		"00000011",	-- 0x394c
		"00000100",	-- 0x394d
		"10111010",	-- 0x394e
		"00000010",	-- 0x394f
		"00010011",	-- 0x3950
		"11111010",	-- 0x3951
		"00000011",	-- 0x3952
		"00000110",	-- 0x3953
		"10110010",	-- 0x3954
		"00000010",	-- 0x3955
		"00010101",	-- 0x3956
		"11111010",	-- 0x3957
		"00000001",	-- 0x3958
		"10111101",	-- 0x3959
		"10110010",	-- 0x395a
		"00000010",	-- 0x395b
		"00011100",	-- 0x395c
		"10010110",	-- 0x395d
		"01001011",	-- 0x395e
		"10111010",	-- 0x395f
		"00000010",	-- 0x3960
		"00011110",	-- 0x3961
		"11011010",	-- 0x3962
		"01000110",	-- 0x3963
		"10110010",	-- 0x3964
		"00000010",	-- 0x3965
		"00100000",	-- 0x3966
		"01010010",	-- 0x3967
		"11111011",	-- 0x3968
		"00000001",	-- 0x3969
		"11010101",	-- 0x396a
		"11001111",	-- 0x396b
		"10000000",	-- 0x396c
		"01000111",	-- 0x396d
		"00000010",	-- 0x396e
		"11000110",	-- 0x396f
		"00000001",	-- 0x3970
		"11111011",	-- 0x3971
		"00000001",	-- 0x3972
		"11011001",	-- 0x3973
		"11001111",	-- 0x3974
		"00000100",	-- 0x3975
		"01000111",	-- 0x3976
		"00000010",	-- 0x3977
		"11000110",	-- 0x3978
		"00000010",	-- 0x3979
		"00110111",	-- 0x397a
		"00111001",	-- 0x397b
		"00000010",	-- 0x397c
		"11000110",	-- 0x397d
		"00000100",	-- 0x397e
		"11111011",	-- 0x397f
		"00000001",	-- 0x3980
		"11010111",	-- 0x3981
		"11001111",	-- 0x3982
		"00000001",	-- 0x3983
		"01000111",	-- 0x3984
		"00000010",	-- 0x3985
		"11000110",	-- 0x3986
		"00001000",	-- 0x3987
		"00110111",	-- 0x3988
		"01011101",	-- 0x3989
		"00000010",	-- 0x398a
		"11000110",	-- 0x398b
		"00010000",	-- 0x398c
		"00110111",	-- 0x398d
		"01111001",	-- 0x398e
		"00000010",	-- 0x398f
		"11000110",	-- 0x3990
		"00100000",	-- 0x3991
		"10110010",	-- 0x3992
		"00000010",	-- 0x3993
		"00100001",	-- 0x3994
		"11011010",	-- 0x3995
		"01000011",	-- 0x3996
		"10110010",	-- 0x3997
		"00000010",	-- 0x3998
		"00100010",	-- 0x3999
		"01100011",	-- 0x399a
		"10001110",	-- 0x399b
		"00000010",	-- 0x399c
		"00100110",	-- 0x399d
		"10001111",	-- 0x399e
		"00000001",	-- 0x399f
		"11011110",	-- 0x39a0
		"00011011",	-- 0x39a1
		"10101010",	-- 0x39a2
		"00000000",	-- 0x39a3
		"00011100",	-- 0x39a4
		"00011100",	-- 0x39a5
		"10001100",	-- 0x39a6
		"00000010",	-- 0x39a7
		"01001000",	-- 0x39a8
		"01000101",	-- 0x39a9
		"11110110",	-- 0x39aa
		"01100011",	-- 0x39ab
		"01110101",	-- 0x39ac
		"00101101",	-- 0x39ad
		"01101110",	-- 0x39ae
		"01101111",	-- 0x39af
		"01110001",	-- 0x39b0
		"01110010",	-- 0x39b1
		"01000110",	-- 0x39b2
		"00000011",	-- 0x39b3
		"00000001",	-- 0x39b4
		"11110000",	-- 0x39b5
		"01011001",	-- 0x39b6
		"01110001",	-- 0x39b7
		"01010010",	-- 0x39b8
		"01000110",	-- 0x39b9
		"00000011",	-- 0x39ba
		"00000001",	-- 0x39bb
		"11110111",	-- 0x39bc
		"11000111",	-- 0x39bd
		"01111111",	-- 0x39be
		"01111110",	-- 0x39bf
		"01110011",	-- 0x39c0
		"01110101",	-- 0x39c1
		"11101101",	-- 0x39c2
		"01101110",	-- 0x39c3
		"01101111",	-- 0x39c4
		"01110001",	-- 0x39c5
		"10100100",	-- 0x39c6
		"01000111",	-- 0x39c7
		"00000101",	-- 0x39c8
		"01110101",	-- 0x39c9
		"10100100",	-- 0x39ca
		"10010110",	-- 0x39cb
		"00011010",	-- 0x39cc
		"10001100",	-- 0x39cd
		"10010110",	-- 0x39ce
		"00110100",	-- 0x39cf
		"01111001",	-- 0x39d0
		"00000101",	-- 0x39d1
		"10110011",	-- 0x39d2
		"01000010",	-- 0x39d3
		"00001001",	-- 0x39d4
		"10011000",	-- 0x39d5
		"01110001",	-- 0x39d6
		"10001001",	-- 0x39d7
		"00000000",	-- 0x39d8
		"11111010",	-- 0x39d9
		"01000011",	-- 0x39da
		"00001111",	-- 0x39db
		"10010111",	-- 0x39dc
		"01110001",	-- 0x39dd
		"10011010",	-- 0x39de
		"01110001",	-- 0x39df
		"00000101",	-- 0x39e0
		"11011010",	-- 0x39e1
		"01101111",	-- 0x39e2
		"01010110",	-- 0x39e3
		"01000111",	-- 0x39e4
		"00000010",	-- 0x39e5
		"10010010",	-- 0x39e6
		"01101111",	-- 0x39e7
		"00000111",	-- 0x39e8
		"01110010",	-- 0x39e9
		"10110011",	-- 0x39ea
		"01000000",	-- 0x39eb
		"00011000",	-- 0x39ec
		"01010010",	-- 0x39ed
		"10001110",	-- 0x39ee
		"00000000",	-- 0x39ef
		"01101111",	-- 0x39f0
		"01101010",	-- 0x39f1
		"00000000",	-- 0x39f2
		"01101010",	-- 0x39f3
		"00000001",	-- 0x39f4
		"11100000",	-- 0x39f5
		"00000001",	-- 0x39f6
		"01000100",	-- 0x39f7
		"00000010",	-- 0x39f8
		"11001010",	-- 0x39f9
		"11111111",	-- 0x39fa
		"11001100",	-- 0x39fb
		"00000010",	-- 0x39fc
		"01000010",	-- 0x39fd
		"00000001",	-- 0x39fe
		"01010010",	-- 0x39ff
		"01111010",	-- 0x3a00
		"01011101",	-- 0x3a01
		"10010010",	-- 0x3a02
		"01110011",	-- 0x3a03
		"01100011",	-- 0x3a04
		"01111111",	-- 0x3a05
		"01111110",	-- 0x3a06
		"01110011",	-- 0x3a07
		"01110101",	-- 0x3a08
		"01101101",	-- 0x3a09
		"01101110",	-- 0x3a0a
		"01101111",	-- 0x3a0b
		"00110101",	-- 0x3a0c
		"11001011",	-- 0x3a0d
		"00001111",	-- 0x3a0e
		"11011010",	-- 0x3a0f
		"00000110",	-- 0x3a10
		"01110111",	-- 0x3a11
		"00101011",	-- 0x3a12
		"00110011",	-- 0x3a13
		"00000010",	-- 0x3a14
		"00000110",	-- 0x3a15
		"11001011",	-- 0x3a16
		"00001101",	-- 0x3a17
		"00110101",	-- 0x3a18
		"11101011",	-- 0x3a19
		"00001001",	-- 0x3a1a
		"01010001",	-- 0x3a1b
		"01000110",	-- 0x3a1c
		"11111010",	-- 0x3a1d
		"11011011",	-- 0x3a1e
		"00000110",	-- 0x3a1f
		"11001010",	-- 0x3a20
		"11111111",	-- 0x3a21
		"01000000",	-- 0x3a22
		"00011101",	-- 0x3a23
		"01110101",	-- 0x3a24
		"01101101",	-- 0x3a25
		"00110101",	-- 0x3a26
		"11001011",	-- 0x3a27
		"11110101",	-- 0x3a28
		"11011011",	-- 0x3a29
		"00000110",	-- 0x3a2a
		"00111110",	-- 0x3a2b
		"00110111",	-- 0x3a2c
		"00110010",	-- 0x3a2d
		"00000011",	-- 0x3a2e
		"00110111",	-- 0x3a2f
		"11110010",	-- 0x3a30
		"00001101",	-- 0x3a31
		"01111001",	-- 0x3a32
		"00011000",	-- 0x3a33
		"10101101",	-- 0x3a34
		"01000010",	-- 0x3a35
		"00001000",	-- 0x3a36
		"01110001",	-- 0x3a37
		"00000000",	-- 0x3a38
		"01000111",	-- 0x3a39
		"00000010",	-- 0x3a3a
		"01110101",	-- 0x3a3b
		"00000000",	-- 0x3a3c
		"01110101",	-- 0x3a3d
		"11110010",	-- 0x3a3e
		"11011010",	-- 0x3a3f
		"11111101",	-- 0x3a40
		"01101100",	-- 0x3a41
		"00110101",	-- 0x3a42
		"00110010",	-- 0x3a43
		"00001101",	-- 0x3a44
		"01010010",	-- 0x3a45
		"11011011",	-- 0x3a46
		"11111101",	-- 0x3a47
		"01010111",	-- 0x3a48
		"11001101",	-- 0x3a49
		"00001110",	-- 0x3a4a
		"01000110",	-- 0x3a4b
		"00110100",	-- 0x3a4c
		"01110111",	-- 0x3a4d
		"00110010",	-- 0x3a4e
		"00000011",	-- 0x3a4f
		"11111010",	-- 0x3a50
		"11001001",	-- 0x3a51
		"11011010",	-- 0x3a52
		"11111110",	-- 0x3a53
		"01010110",	-- 0x3a54
		"11000010",	-- 0x3a55
		"01111111",	-- 0x3a56
		"01011011",	-- 0x3a57
		"11000011",	-- 0x3a58
		"00000111",	-- 0x3a59
		"10001111",	-- 0x3a5a
		"11111010",	-- 0x3a5b
		"11111010",	-- 0x3a5c
		"00110101",	-- 0x3a5d
		"00110000",	-- 0x3a5e
		"00000110",	-- 0x3a5f
		"00110101",	-- 0x3a60
		"00010000",	-- 0x3a61
		"00000011",	-- 0x3a62
		"10001111",	-- 0x3a63
		"11111011",	-- 0x3a64
		"00000010",	-- 0x3a65
		"00001111",	-- 0x3a66
		"11101011",	-- 0x3a67
		"10000000",	-- 0x3a68
		"01001010",	-- 0x3a69
		"00010110",	-- 0x3a6a
		"11001101",	-- 0x3a6b
		"10000001",	-- 0x3a6c
		"01000111",	-- 0x3a6d
		"00000110",	-- 0x3a6e
		"11001101",	-- 0x3a6f
		"10000000",	-- 0x3a70
		"01000111",	-- 0x3a71
		"00011010",	-- 0x3a72
		"01000000",	-- 0x3a73
		"01010010",	-- 0x3a74
		"01011011",	-- 0x3a75
		"00010001",	-- 0x3a76
		"00010001",	-- 0x3a77
		"00010001",	-- 0x3a78
		"11000011",	-- 0x3a79
		"00001111",	-- 0x3a7a
		"10001111",	-- 0x3a7b
		"11111011",	-- 0x3a7c
		"00001010",	-- 0x3a7d
		"00001111",	-- 0x3a7e
		"11101011",	-- 0x3a7f
		"10000000",	-- 0x3a80
		"01110111",	-- 0x3a81
		"00101011",	-- 0x3a82
		"10010011",	-- 0x3a83
		"11111101",	-- 0x3a84
		"01100111",	-- 0x3a85
		"00010111",	-- 0x3a86
		"11000011",	-- 0x3a87
		"00011111",	-- 0x3a88
		"10010011",	-- 0x3a89
		"00000110",	-- 0x3a8a
		"01000000",	-- 0x3a8b
		"00111010",	-- 0x3a8c
		"01101100",	-- 0x3a8d
		"01110101",	-- 0x3a8e
		"00101011",	-- 0x3a8f
		"11001010",	-- 0x3a90
		"11011010",	-- 0x3a91
		"10010010",	-- 0x3a92
		"00000110",	-- 0x3a93
		"11001010",	-- 0x3a94
		"00001110",	-- 0x3a95
		"00110101",	-- 0x3a96
		"11101011",	-- 0x3a97
		"00000101",	-- 0x3a98
		"01010000",	-- 0x3a99
		"01000110",	-- 0x3a9a
		"11111010",	-- 0x3a9b
		"01000000",	-- 0x3a9c
		"00000011",	-- 0x3a9d
		"00110111",	-- 0x3a9e
		"11001011",	-- 0x3a9f
		"00000100",	-- 0x3aa0
		"11011010",	-- 0x3aa1
		"00000110",	-- 0x3aa2
		"01000000",	-- 0x3aa3
		"00011100",	-- 0x3aa4
		"11011011",	-- 0x3aa5
		"00000110",	-- 0x3aa6
		"11011010",	-- 0x3aa7
		"00101011",	-- 0x3aa8
		"11000010",	-- 0x3aa9
		"00000001",	-- 0x3aaa
		"10001001",	-- 0x3aab
		"00000000",	-- 0x3aac
		"00011111",	-- 0x3aad
		"01000110",	-- 0x3aae
		"00000100",	-- 0x3aaf
		"10000110",	-- 0x3ab0
		"11111111",	-- 0x3ab1
		"11011100",	-- 0x3ab2
		"01000001",	-- 0x3ab3
		"00000110",	-- 0x3ab4
		"00111111",	-- 0x3ab5
		"00011011",	-- 0x3ab6
		"01110101",	-- 0x3ab7
		"00101011",	-- 0x3ab8
		"10010010",	-- 0x3ab9
		"00000110",	-- 0x3aba
		"10000101",	-- 0x3abb
		"00000000",	-- 0x3abc
		"01110101",	-- 0x3abd
		"00101011",	-- 0x3abe
		"10010011",	-- 0x3abf
		"00000110",	-- 0x3ac0
		"01110101",	-- 0x3ac1
		"01101101",	-- 0x3ac2
		"01111100",	-- 0x3ac3
		"01010110",	-- 0x3ac4
		"11000010",	-- 0x3ac5
		"01111111",	-- 0x3ac6
		"10010010",	-- 0x3ac7
		"11111110",	-- 0x3ac8
		"01111101",	-- 0x3ac9
		"11001101",	-- 0x3aca
		"11111111",	-- 0x3acb
		"01000110",	-- 0x3acc
		"00000011",	-- 0x3acd
		"00000011",	-- 0x3ace
		"11111011",	-- 0x3acf
		"00011010",	-- 0x3ad0
		"00010011",	-- 0x3ad1
		"11000011",	-- 0x3ad2
		"00011110",	-- 0x3ad3
		"10001111",	-- 0x3ad4
		"11111010",	-- 0x3ad5
		"11011110",	-- 0x3ad6
		"00001111",	-- 0x3ad7
		"10101111",	-- 0x3ad8
		"10000000",	-- 0x3ad9
		"00111100",	-- 0x3ada
		"01011011",	-- 0x3adb
		"00100011",	-- 0x3adc
		"10000000",	-- 0x3add
		"11111011",	-- 0x3ade
		"10001010",	-- 0x3adf
		"11111100",	-- 0x3ae0
		"10011011",	-- 0x3ae1
		"11111100",	-- 0x3ae2
		"01011101",	-- 0x3ae3
		"11111111",	-- 0x3ae4
		"01011000",	-- 0x3ae5
		"11111111",	-- 0x3ae6
		"01111011",	-- 0x3ae7
		"11111110",	-- 0x3ae8
		"11101010",	-- 0x3ae9
		"11111111",	-- 0x3aea
		"10111110",	-- 0x3aeb
		"11111111",	-- 0x3aec
		"11000100",	-- 0x3aed
		"11111110",	-- 0x3aee
		"00010101",	-- 0x3aef
		"11111111",	-- 0x3af0
		"11001010",	-- 0x3af1
		"11111111",	-- 0x3af2
		"00100001",	-- 0x3af3
		"11111111",	-- 0x3af4
		"11010110",	-- 0x3af5
		"11111111",	-- 0x3af6
		"10111000",	-- 0x3af7
		"11111111",	-- 0x3af8
		"11010000",	-- 0x3af9
		"10000010",	-- 0x3afa
		"00000010",	-- 0x3afb
		"10000001",	-- 0x3afc
		"10000000",	-- 0x3afd
		"10000010",	-- 0x3afe
		"00001000",	-- 0x3aff
		"00000001",	-- 0x3b00
		"10000000",	-- 0x3b01
		"10000010",	-- 0x3b02
		"00000011",	-- 0x3b03
		"10000001",	-- 0x3b04
		"10000000",	-- 0x3b05
		"10000010",	-- 0x3b06
		"00001000",	-- 0x3b07
		"00000001",	-- 0x3b08
		"10000000",	-- 0x3b09
		"00000100",	-- 0x3b0a
		"00001010",	-- 0x3b0b
		"00000011",	-- 0x3b0c
		"00000110",	-- 0x3b0d
		"00000100",	-- 0x3b0e
		"00000101",	-- 0x3b0f
		"00000011",	-- 0x3b10
		"00000111",	-- 0x3b11
		"00000100",	-- 0x3b12
		"00001010",	-- 0x3b13
		"00000011",	-- 0x3b14
		"00001001",	-- 0x3b15
		"00000100",	-- 0x3b16
		"00001101",	-- 0x3b17
		"00000011",	-- 0x3b18
		"00001100",	-- 0x3b19
		"01111111",	-- 0x3b1a
		"01111110",	-- 0x3b1b
		"01110011",	-- 0x3b1c
		"01010010",	-- 0x3b1d
		"00110111",	-- 0x3b1e
		"00100000",	-- 0x3b1f
		"00000010",	-- 0x3b20
		"11000110",	-- 0x3b21
		"00000001",	-- 0x3b22
		"00110101",	-- 0x3b23
		"01000000",	-- 0x3b24
		"00000010",	-- 0x3b25
		"11000110",	-- 0x3b26
		"00000010",	-- 0x3b27
		"00110101",	-- 0x3b28
		"01100000",	-- 0x3b29
		"00000010",	-- 0x3b2a
		"11000110",	-- 0x3b2b
		"00000100",	-- 0x3b2c
		"00110101",	-- 0x3b2d
		"10000000",	-- 0x3b2e
		"00000010",	-- 0x3b2f
		"11000110",	-- 0x3b30
		"00001000",	-- 0x3b31
		"00110111",	-- 0x3b32
		"10100000",	-- 0x3b33
		"00000010",	-- 0x3b34
		"11000110",	-- 0x3b35
		"00010000",	-- 0x3b36
		"00110101",	-- 0x3b37
		"11000010",	-- 0x3b38
		"00000010",	-- 0x3b39
		"11000110",	-- 0x3b3a
		"00100000",	-- 0x3b3b
		"00110101",	-- 0x3b3c
		"11100010",	-- 0x3b3d
		"00000010",	-- 0x3b3e
		"11000110",	-- 0x3b3f
		"01000000",	-- 0x3b40
		"00110111",	-- 0x3b41
		"01001001",	-- 0x3b42
		"00000010",	-- 0x3b43
		"11000110",	-- 0x3b44
		"10000000",	-- 0x3b45
		"10001110",	-- 0x3b46
		"00000000",	-- 0x3b47
		"01001001",	-- 0x3b48
		"10001111",	-- 0x3b49
		"00000001",	-- 0x3b4a
		"00000011",	-- 0x3b4b
		"01100001",	-- 0x3b4c
		"00101111",	-- 0x3b4d
		"01010010",	-- 0x3b4e
		"00110111",	-- 0x3b4f
		"01101001",	-- 0x3b50
		"00000010",	-- 0x3b51
		"11000110",	-- 0x3b52
		"00000001",	-- 0x3b53
		"00110111",	-- 0x3b54
		"00001000",	-- 0x3b55
		"00000010",	-- 0x3b56
		"11000110",	-- 0x3b57
		"00000010",	-- 0x3b58
		"00110101",	-- 0x3b59
		"00101000",	-- 0x3b5a
		"00000010",	-- 0x3b5b
		"11000110",	-- 0x3b5c
		"00000100",	-- 0x3b5d
		"00110101",	-- 0x3b5e
		"01001000",	-- 0x3b5f
		"00000010",	-- 0x3b60
		"11000110",	-- 0x3b61
		"00001000",	-- 0x3b62
		"00110101",	-- 0x3b63
		"11001000",	-- 0x3b64
		"00000010",	-- 0x3b65
		"11000110",	-- 0x3b66
		"00010000",	-- 0x3b67
		"00110101",	-- 0x3b68
		"11101000",	-- 0x3b69
		"00000010",	-- 0x3b6a
		"11000110",	-- 0x3b6b
		"00100000",	-- 0x3b6c
		"00110101",	-- 0x3b6d
		"00001101",	-- 0x3b6e
		"00000010",	-- 0x3b6f
		"11000110",	-- 0x3b70
		"01000000",	-- 0x3b71
		"00110111",	-- 0x3b72
		"10000011",	-- 0x3b73
		"00000010",	-- 0x3b74
		"11000110",	-- 0x3b75
		"10000000",	-- 0x3b76
		"10001110",	-- 0x3b77
		"00000000",	-- 0x3b78
		"01001010",	-- 0x3b79
		"10001111",	-- 0x3b7a
		"00000001",	-- 0x3b7b
		"00000100",	-- 0x3b7c
		"01011011",	-- 0x3b7d
		"11101000",	-- 0x3b7e
		"00000000",	-- 0x3b7f
		"11100010",	-- 0x3b80
		"10000000",	-- 0x3b81
		"10100011",	-- 0x3b82
		"10000000",	-- 0x3b83
		"11100011",	-- 0x3b84
		"00000000",	-- 0x3b85
		"00001000",	-- 0x3b86
		"10100010",	-- 0x3b87
		"00000000",	-- 0x3b88
		"01100011",	-- 0x3b89
		"10001111",	-- 0x3b8a
		"11000011",	-- 0x3b8b
		"11000111",	-- 0x3b8c
		"00100001",	-- 0x3b8d
		"10010000",	-- 0x3b8e
		"11111010",	-- 0x3b8f
		"00000001",	-- 0x3b90
		"10001100",	-- 0x3b91
		"01000100",	-- 0x3b92
		"00100010",	-- 0x3b93
		"10001110",	-- 0x3b94
		"01100110",	-- 0x3b95
		"01100110",	-- 0x3b96
		"00110111",	-- 0x3b97
		"01010000",	-- 0x3b98
		"00000100",	-- 0x3b99
		"01110111",	-- 0x3b9a
		"10111011",	-- 0x3b9b
		"01110111",	-- 0x3b9c
		"01111000",	-- 0x3b9d
		"11001110",	-- 0x3b9e
		"00000001",	-- 0x3b9f
		"01000110",	-- 0x3ba0
		"00000110",	-- 0x3ba1
		"11000110",	-- 0x3ba2
		"00000001",	-- 0x3ba3
		"01110010",	-- 0x3ba4
		"11011111",	-- 0x3ba5
		"01000000",	-- 0x3ba6
		"00010111",	-- 0x3ba7
		"01111001",	-- 0x3ba8
		"00001111",	-- 0x3ba9
		"11011111",	-- 0x3baa
		"01000101",	-- 0x3bab
		"00000010",	-- 0x3bac
		"01110111",	-- 0x3bad
		"10111011",	-- 0x3bae
		"10001110",	-- 0x3baf
		"01100110",	-- 0x3bb0
		"01100110",	-- 0x3bb1
		"01110111",	-- 0x3bb2
		"01111101",	-- 0x3bb3
		"01000000",	-- 0x3bb4
		"00001001",	-- 0x3bb5
		"11000010",	-- 0x3bb6
		"11111110",	-- 0x3bb7
		"00110101",	-- 0x3bb8
		"01010000",	-- 0x3bb9
		"00000010",	-- 0x3bba
		"01110101",	-- 0x3bbb
		"10111011",	-- 0x3bbc
		"01110101",	-- 0x3bbd
		"01111101",	-- 0x3bbe
		"10110010",	-- 0x3bbf
		"00000001",	-- 0x3bc0
		"10001100",	-- 0x3bc1
		"00111100",	-- 0x3bc2
		"10001000",	-- 0x3bc3
		"00101001",	-- 0x3bc4
		"01000000",	-- 0x3bc5
		"01000100",	-- 0x3bc6
		"00000100",	-- 0x3bc7
		"01010010",	-- 0x3bc8
		"01010011",	-- 0x3bc9
		"01000000",	-- 0x3bca
		"00010100",	-- 0x3bcb
		"00111110",	-- 0x3bcc
		"01101101",	-- 0x3bcd
		"10000001",	-- 0x3bce
		"01001001",	-- 0x3bcf
		"10111010",	-- 0x3bd0
		"00000001",	-- 0x3bd1
		"00100101",	-- 0x3bd2
		"01111100",	-- 0x3bd3
		"10000001",	-- 0x3bd4
		"01001001",	-- 0x3bd5
		"00001100",	-- 0x3bd6
		"00111100",	-- 0x3bd7
		"10110111",	-- 0x3bd8
		"00000001",	-- 0x3bd9
		"00100101",	-- 0x3bda
		"01000100",	-- 0x3bdb
		"00000011",	-- 0x3bdc
		"10000110",	-- 0x3bdd
		"11111111",	-- 0x3bde
		"11111111",	-- 0x3bdf
		"00110101",	-- 0x3be0
		"00010000",	-- 0x3be1
		"01001101",	-- 0x3be2
		"00110101",	-- 0x3be3
		"00110111",	-- 0x3be4
		"00010000",	-- 0x3be5
		"01111001",	-- 0x3be6
		"00001100",	-- 0x3be7
		"00000100",	-- 0x3be8
		"01000101",	-- 0x3be9
		"01000101",	-- 0x3bea
		"01110111",	-- 0x3beb
		"00110111",	-- 0x3bec
		"10010010",	-- 0x3bed
		"11111010",	-- 0x3bee
		"00110111",	-- 0x3bef
		"00011001",	-- 0x3bf0
		"00111110",	-- 0x3bf1
		"01110111",	-- 0x3bf2
		"01010111",	-- 0x3bf3
		"01000000",	-- 0x3bf4
		"00111010",	-- 0x3bf5
		"10011000",	-- 0x3bf6
		"01010000",	-- 0x3bf7
		"00010100",	-- 0x3bf8
		"00010101",	-- 0x3bf9
		"00000001",	-- 0x3bfa
		"11000100",	-- 0x3bfb
		"11010111",	-- 0x3bfc
		"10010111",	-- 0x3bfd
		"01010000",	-- 0x3bfe
		"00111111",	-- 0x3bff
		"00110101",	-- 0x3c00
		"01010111",	-- 0x3c01
		"00010110",	-- 0x3c02
		"11010100",	-- 0x3c03
		"11111010",	-- 0x3c04
		"01000100",	-- 0x3c05
		"00000001",	-- 0x3c06
		"01010100",	-- 0x3c07
		"11001100",	-- 0x3c08
		"00000001",	-- 0x3c09
		"00111101",	-- 0x3c0a
		"01000010",	-- 0x3c0b
		"11100101",	-- 0x3c0c
		"00110111",	-- 0x3c0d
		"00011001",	-- 0x3c0e
		"00001001",	-- 0x3c0f
		"01110111",	-- 0x3c10
		"01010111",	-- 0x3c11
		"01111001",	-- 0x3c12
		"11111111",	-- 0x3c13
		"11000111",	-- 0x3c14
		"01000101",	-- 0x3c15
		"00000010",	-- 0x3c16
		"01110111",	-- 0x3c17
		"00010111",	-- 0x3c18
		"00110111",	-- 0x3c19
		"00010111",	-- 0x3c1a
		"00010100",	-- 0x3c1b
		"00110111",	-- 0x3c1c
		"10101010",	-- 0x3c1d
		"00010001",	-- 0x3c1e
		"01101000",	-- 0x3c1f
		"11011011",	-- 0x3c20
		"11111010",	-- 0x3c21
		"10001111",	-- 0x3c22
		"11000011",	-- 0x3c23
		"10111101",	-- 0x3c24
		"00100001",	-- 0x3c25
		"10011010",	-- 0x3c26
		"10001110",	-- 0x3c27
		"00000000",	-- 0x3c28
		"10011000",	-- 0x3c29
		"00000001",	-- 0x3c2a
		"11010001",	-- 0x3c2b
		"10011000",	-- 0x3c2c
		"01110101",	-- 0x3c2d
		"00010111",	-- 0x3c2e
		"01111000",	-- 0x3c2f
		"10011010",	-- 0x3c30
		"01010000",	-- 0x3c31
		"10111010",	-- 0x3c32
		"00000010",	-- 0x3c33
		"00000000",	-- 0x3c34
		"00000011",	-- 0x3c35
		"11111100",	-- 0x3c36
		"01010111",	-- 0x3c37
		"11011011",	-- 0x3c38
		"10011000",	-- 0x3c39
		"10001111",	-- 0x3c3a
		"11000011",	-- 0x3c3b
		"10111101",	-- 0x3c3c
		"00100001",	-- 0x3c3d
		"10011010",	-- 0x3c3e
		"01000100",	-- 0x3c3f
		"00000011",	-- 0x3c40
		"00000001",	-- 0x3c41
		"11001000",	-- 0x3c42
		"00001000",	-- 0x3c43
		"11011010",	-- 0x3c44
		"10011000",	-- 0x3c45
		"00110101",	-- 0x3c46
		"00010010",	-- 0x3c47
		"00000010",	-- 0x3c48
		"11001010",	-- 0x3c49
		"01010000",	-- 0x3c4a
		"01010011",	-- 0x3c4b
		"00000100",	-- 0x3c4c
		"10000101",	-- 0x3c4d
		"01100001",	-- 0x3c4e
		"01000100",	-- 0x3c4f
		"00000010",	-- 0x3c50
		"11001011",	-- 0x3c51
		"11111111",	-- 0x3c52
		"10110011",	-- 0x3c53
		"00000001",	-- 0x3c54
		"01000100",	-- 0x3c55
		"01100011",	-- 0x3c56
		"00000001",	-- 0x3c57
		"11001100",	-- 0x3c58
		"11010110",	-- 0x3c59
		"00000011",	-- 0x3c5a
		"11111011",	-- 0x3c5b
		"00011010",	-- 0x3c5c
		"00111100",	-- 0x3c5d
		"00000110",	-- 0x3c5e
		"01000101",	-- 0x3c5f
		"00000011",	-- 0x3c60
		"00000110",	-- 0x3c61
		"01000100",	-- 0x3c62
		"00000010",	-- 0x3c63
		"11001010",	-- 0x3c64
		"11111111",	-- 0x3c65
		"10110010",	-- 0x3c66
		"00000001",	-- 0x3c67
		"10000110",	-- 0x3c68
		"11011011",	-- 0x3c69
		"01011111",	-- 0x3c6a
		"10001111",	-- 0x3c6b
		"11000010",	-- 0x3c6c
		"01001001",	-- 0x3c6d
		"00110101",	-- 0x3c6e
		"01010110",	-- 0x3c6f
		"00001010",	-- 0x3c70
		"00011101",	-- 0x3c71
		"11111010",	-- 0x3c72
		"00000001",	-- 0x3c73
		"00000010",	-- 0x3c74
		"00010010",	-- 0x3c75
		"00010110",	-- 0x3c76
		"00010110",	-- 0x3c77
		"11000010",	-- 0x3c78
		"00000011",	-- 0x3c79
		"00001101",	-- 0x3c7a
		"10001100",	-- 0x3c7b
		"00010111",	-- 0x3c7c
		"00001010",	-- 0x3c7d
		"01000101",	-- 0x3c7e
		"00001001",	-- 0x3c7f
		"11101010",	-- 0x3c80
		"10000101",	-- 0x3c81
		"01010001",	-- 0x3c82
		"01001011",	-- 0x3c83
		"00001101",	-- 0x3c84
		"01000111",	-- 0x3c85
		"00001001",	-- 0x3c86
		"01000000",	-- 0x3c87
		"00001010",	-- 0x3c88
		"11101010",	-- 0x3c89
		"10000000",	-- 0x3c8a
		"01010111",	-- 0x3c8b
		"01001011",	-- 0x3c8c
		"00000101",	-- 0x3c8d
		"01000110",	-- 0x3c8e
		"00000010",	-- 0x3c8f
		"01110111",	-- 0x3c90
		"10010100",	-- 0x3c91
		"01011011",	-- 0x3c92
		"10010011",	-- 0x3c93
		"01011111",	-- 0x3c94
		"10110011",	-- 0x3c95
		"00000010",	-- 0x3c96
		"00010010",	-- 0x3c97
		"00000011",	-- 0x3c98
		"11111011",	-- 0x3c99
		"00011010",	-- 0x3c9a
		"10110011",	-- 0x3c9b
		"00000001",	-- 0x3c9c
		"01001111",	-- 0x3c9d
		"11111010",	-- 0x3c9e
		"00000001",	-- 0x3c9f
		"10001100",	-- 0x3ca0
		"11001101",	-- 0x3ca1
		"00001101",	-- 0x3ca2
		"01000101",	-- 0x3ca3
		"00101000",	-- 0x3ca4
		"11001101",	-- 0x3ca5
		"11111011",	-- 0x3ca6
		"01000010",	-- 0x3ca7
		"00100111",	-- 0x3ca8
		"00110101",	-- 0x3ca9
		"00111001",	-- 0x3caa
		"00000101",	-- 0x3cab
		"00110111",	-- 0x3cac
		"00111100",	-- 0x3cad
		"00001111",	-- 0x3cae
		"01000000",	-- 0x3caf
		"00010110",	-- 0x3cb0
		"11001101",	-- 0x3cb1
		"01001101",	-- 0x3cb2
		"01000100",	-- 0x3cb3
		"00011011",	-- 0x3cb4
		"11001101",	-- 0x3cb5
		"00110001",	-- 0x3cb6
		"01000010",	-- 0x3cb7
		"00001110",	-- 0x3cb8
		"00110101",	-- 0x3cb9
		"01010000",	-- 0x3cba
		"00000010",	-- 0x3cbb
		"01110101",	-- 0x3cbc
		"00111100",	-- 0x3cbd
		"11001110",	-- 0x3cbe
		"00100000",	-- 0x3cbf
		"01000111",	-- 0x3cc0
		"00000010",	-- 0x3cc1
		"01110101",	-- 0x3cc2
		"11110000",	-- 0x3cc3
		"11000110",	-- 0x3cc4
		"00100000",	-- 0x3cc5
		"10001100",	-- 0x3cc6
		"11000010",	-- 0x3cc7
		"11011111",	-- 0x3cc8
		"11000010",	-- 0x3cc9
		"11110111",	-- 0x3cca
		"01000000",	-- 0x3ccb
		"00100011",	-- 0x3ccc
		"00110101",	-- 0x3ccd
		"00111001",	-- 0x3cce
		"11110111",	-- 0x3ccf
		"01110111",	-- 0x3cd0
		"11110000",	-- 0x3cd1
		"01110101",	-- 0x3cd2
		"01110110",	-- 0x3cd3
		"11001011",	-- 0x3cd4
		"00010000",	-- 0x3cd5
		"10110011",	-- 0x3cd6
		"00000001",	-- 0x3cd7
		"00000001",	-- 0x3cd8
		"11000010",	-- 0x3cd9
		"11011111",	-- 0x3cda
		"11001110",	-- 0x3cdb
		"00001000",	-- 0x3cdc
		"01000110",	-- 0x3cdd
		"00000100",	-- 0x3cde
		"01110010",	-- 0x3cdf
		"11011111",	-- 0x3ce0
		"11000110",	-- 0x3ce1
		"00001000",	-- 0x3ce2
		"00110101",	-- 0x3ce3
		"01010000",	-- 0x3ce4
		"00000110",	-- 0x3ce5
		"01111001",	-- 0x3ce6
		"00001111",	-- 0x3ce7
		"11011111",	-- 0x3ce8
		"01000101",	-- 0x3ce9
		"00000101",	-- 0x3cea
		"10001100",	-- 0x3ceb
		"01110111",	-- 0x3cec
		"01111000",	-- 0x3ced
		"01110111",	-- 0x3cee
		"00111100",	-- 0x3cef
		"10110010",	-- 0x3cf0
		"00000001",	-- 0x3cf1
		"10001100",	-- 0x3cf2
		"00110111",	-- 0x3cf3
		"11110000",	-- 0x3cf4
		"00001101",	-- 0x3cf5
		"01110010",	-- 0x3cf6
		"11101111",	-- 0x3cf7
		"10000110",	-- 0x3cf8
		"00000000",	-- 0x3cf9
		"00000000",	-- 0x3cfa
		"10011010",	-- 0x3cfb
		"01010010",	-- 0x3cfc
		"10111010",	-- 0x3cfd
		"00000010",	-- 0x3cfe
		"00000010",	-- 0x3cff
		"00000011",	-- 0x3d00
		"11111101",	-- 0x3d01
		"10011110",	-- 0x3d02
		"00110101",	-- 0x3d03
		"00111001",	-- 0x3d04
		"00000010",	-- 0x3d05
		"01110010",	-- 0x3d06
		"11101111",	-- 0x3d07
		"11111010",	-- 0x3d08
		"00000011",	-- 0x3d09
		"00000000",	-- 0x3d0a
		"11001011",	-- 0x3d0b
		"10101110",	-- 0x3d0c
		"00110101",	-- 0x3d0d
		"00010000",	-- 0x3d0e
		"01010111",	-- 0x3d0f
		"00110111",	-- 0x3d10
		"00110010",	-- 0x3d11
		"01010100",	-- 0x3d12
		"00110111",	-- 0x3d13
		"00010010",	-- 0x3d14
		"01010001",	-- 0x3d15
		"01110001",	-- 0x3d16
		"10110111",	-- 0x3d17
		"01000110",	-- 0x3d18
		"00001000",	-- 0x3d19
		"11000000",	-- 0x3d1a
		"00001000",	-- 0x3d1b
		"01000100",	-- 0x3d1c
		"00000010",	-- 0x3d1d
		"11001010",	-- 0x3d1e
		"11111111",	-- 0x3d1f
		"01000000",	-- 0x3d20
		"00110101",	-- 0x3d21
		"11011011",	-- 0x3d22
		"11101111",	-- 0x3d23
		"11001101",	-- 0x3d24
		"01000000",	-- 0x3d25
		"01000101",	-- 0x3d26
		"00000100",	-- 0x3d27
		"11000101",	-- 0x3d28
		"01000000",	-- 0x3d29
		"01000000",	-- 0x3d2a
		"11111000",	-- 0x3d2b
		"11001101",	-- 0x3d2c
		"00001010",	-- 0x3d2d
		"01000110",	-- 0x3d2e
		"00001010",	-- 0x3d2f
		"11000000",	-- 0x3d30
		"00000001",	-- 0x3d31
		"01000100",	-- 0x3d32
		"00000010",	-- 0x3d33
		"11001010",	-- 0x3d34
		"11111111",	-- 0x3d35
		"01110110",	-- 0x3d36
		"11101111",	-- 0x3d37
		"01000000",	-- 0x3d38
		"00011101",	-- 0x3d39
		"01111001",	-- 0x3d3a
		"00000010",	-- 0x3d3b
		"11101111",	-- 0x3d3c
		"01000101",	-- 0x3d3d
		"00101001",	-- 0x3d3e
		"01101100",	-- 0x3d3f
		"00111100",	-- 0x3d40
		"00000001",	-- 0x3d41
		"11000100",	-- 0x3d42
		"11011011",	-- 0x3d43
		"11000001",	-- 0x3d44
		"00000001",	-- 0x3d45
		"01000100",	-- 0x3d46
		"00000010",	-- 0x3d47
		"11001011",	-- 0x3d48
		"11111111",	-- 0x3d49
		"01111100",	-- 0x3d4a
		"00001011",	-- 0x3d4b
		"01000011",	-- 0x3d4c
		"00011010",	-- 0x3d4d
		"01110001",	-- 0x3d4e
		"10110010",	-- 0x3d4f
		"01000111",	-- 0x3d50
		"00011000",	-- 0x3d51
		"11000100",	-- 0x3d52
		"00000001",	-- 0x3d53
		"01000100",	-- 0x3d54
		"00000001",	-- 0x3d55
		"01010010",	-- 0x3d56
		"01011011",	-- 0x3d57
		"10001111",	-- 0x3d58
		"11000011",	-- 0x3d59
		"11010011",	-- 0x3d5a
		"00100001",	-- 0x3d5b
		"10000100",	-- 0x3d5c
		"01101110",	-- 0x3d5d
		"10001110",	-- 0x3d5e
		"00000011",	-- 0x3d5f
		"00000000",	-- 0x3d60
		"00000001",	-- 0x3d61
		"11010001",	-- 0x3d62
		"10011000",	-- 0x3d63
		"01111110",	-- 0x3d64
		"01000000",	-- 0x3d65
		"00000011",	-- 0x3d66
		"01011010",	-- 0x3d67
		"01110101",	-- 0x3d68
		"10110010",	-- 0x3d69
		"01010011",	-- 0x3d6a
		"00000100",	-- 0x3d6b
		"00000100",	-- 0x3d6c
		"01101000",	-- 0x3d6d
		"00111100",	-- 0x3d6e
		"00101110",	-- 0x3d6f
		"10101000",	-- 0x3d70
		"00000000",	-- 0x3d71
		"01000100",	-- 0x3d72
		"00000010",	-- 0x3d73
		"01010010",	-- 0x3d74
		"01010011",	-- 0x3d75
		"10111010",	-- 0x3d76
		"00000001",	-- 0x3d77
		"01010000",	-- 0x3d78
		"01111110",	-- 0x3d79
		"10110110",	-- 0x3d7a
		"00000001",	-- 0x3d7b
		"01010010",	-- 0x3d7c
		"10000111",	-- 0x3d7d
		"00000011",	-- 0x3d7e
		"01111011",	-- 0x3d7f
		"01000101",	-- 0x3d80
		"00000101",	-- 0x3d81
		"10111001",	-- 0x3d82
		"00000001",	-- 0x3d83
		"01010000",	-- 0x3d84
		"01000011",	-- 0x3d85
		"00000011",	-- 0x3d86
		"10110110",	-- 0x3d87
		"00000001",	-- 0x3d88
		"01010000",	-- 0x3d89
		"10011010",	-- 0x3d8a
		"01010010",	-- 0x3d8b
		"10111010",	-- 0x3d8c
		"00000010",	-- 0x3d8d
		"00000010",	-- 0x3d8e
		"11001011",	-- 0x3d8f
		"01001100",	-- 0x3d90
		"00110101",	-- 0x3d91
		"01110110",	-- 0x3d92
		"00000010",	-- 0x3d93
		"11001011",	-- 0x3d94
		"01010010",	-- 0x3d95
		"00001011",	-- 0x3d96
		"01000101",	-- 0x3d97
		"00000011",	-- 0x3d98
		"01110111",	-- 0x3d99
		"01110110",	-- 0x3d9a
		"10001100",	-- 0x3d9b
		"01110101",	-- 0x3d9c
		"01110110",	-- 0x3d9d
		"00110111",	-- 0x3d9e
		"11110000",	-- 0x3d9f
		"00001001",	-- 0x3da0
		"01010010",	-- 0x3da1
		"10010010",	-- 0x3da2
		"01011110",	-- 0x3da3
		"01110101",	-- 0x3da4
		"11010111",	-- 0x3da5
		"01110111",	-- 0x3da6
		"11110111",	-- 0x3da7
		"01000000",	-- 0x3da8
		"01011011",	-- 0x3da9
		"10011110",	-- 0x3daa
		"11111111",	-- 0x3dab
		"10010110",	-- 0x3dac
		"01010010",	-- 0x3dad
		"01101110",	-- 0x3dae
		"00101110",	-- 0x3daf
		"10101000",	-- 0x3db0
		"00000000",	-- 0x3db1
		"01111110",	-- 0x3db2
		"01000100",	-- 0x3db3
		"00010111",	-- 0x3db4
		"01010100",	-- 0x3db5
		"01010101",	-- 0x3db6
		"10000100",	-- 0x3db7
		"00000000",	-- 0x3db8
		"10001001",	-- 0x3db9
		"00111101",	-- 0x3dba
		"01110001",	-- 0x3dbb
		"01000101",	-- 0x3dbc
		"00000010",	-- 0x3dbd
		"01110111",	-- 0x3dbe
		"11110111",	-- 0x3dbf
		"11001110",	-- 0x3dc0
		"11100000",	-- 0x3dc1
		"01000110",	-- 0x3dc2
		"00000100",	-- 0x3dc3
		"00000110",	-- 0x3dc4
		"00000110",	-- 0x3dc5
		"01010100",	-- 0x3dc6
		"10001100",	-- 0x3dc7
		"11001010",	-- 0x3dc8
		"10000000",	-- 0x3dc9
		"01000000",	-- 0x3dca
		"00001111",	-- 0x3dcb
		"11001100",	-- 0x3dcc
		"00110011",	-- 0x3dcd
		"01000101",	-- 0x3dce
		"00000010",	-- 0x3dcf
		"01110111",	-- 0x3dd0
		"10110011",	-- 0x3dd1
		"11001110",	-- 0x3dd2
		"11100000",	-- 0x3dd3
		"01000110",	-- 0x3dd4
		"00000011",	-- 0x3dd5
		"00000110",	-- 0x3dd6
		"00000110",	-- 0x3dd7
		"10001100",	-- 0x3dd8
		"11001010",	-- 0x3dd9
		"01111111",	-- 0x3dda
		"11111011",	-- 0x3ddb
		"00000001",	-- 0x3ddc
		"01000110",	-- 0x3ddd
		"01001010",	-- 0x3dde
		"00000001",	-- 0x3ddf
		"01010101",	-- 0x3de0
		"11001101",	-- 0x3de1
		"00000001",	-- 0x3de2
		"01000100",	-- 0x3de3
		"00000010",	-- 0x3de4
		"01110101",	-- 0x3de5
		"11110111",	-- 0x3de6
		"11011011",	-- 0x3de7
		"01011110",	-- 0x3de8
		"10010010",	-- 0x3de9
		"01011110",	-- 0x3dea
		"00110101",	-- 0x3deb
		"01010110",	-- 0x3dec
		"00010101",	-- 0x3ded
		"01111001",	-- 0x3dee
		"10100000",	-- 0x3def
		"01011011",	-- 0x3df0
		"01000100",	-- 0x3df1
		"00010000",	-- 0x3df2
		"00001000",	-- 0x3df3
		"01001001",	-- 0x3df4
		"00001010",	-- 0x3df5
		"01011000",	-- 0x3df6
		"01000111",	-- 0x3df7
		"00001010",	-- 0x3df8
		"01001010",	-- 0x3df9
		"00000001",	-- 0x3dfa
		"01010100",	-- 0x3dfb
		"11001100",	-- 0x3dfc
		"00000010",	-- 0x3dfd
		"01000101",	-- 0x3dfe
		"00000101",	-- 0x3dff
		"01110111",	-- 0x3e00
		"11010111",	-- 0x3e01
		"10001100",	-- 0x3e02
		"01110101",	-- 0x3e03
		"11010111",	-- 0x3e04
		"10010110",	-- 0x3e05
		"01010010",	-- 0x3e06
		"10011010",	-- 0x3e07
		"11111111",	-- 0x3e08
		"00000001",	-- 0x3e09
		"11001001",	-- 0x3e0a
		"10010110",	-- 0x3e0b
		"00000001",	-- 0x3e0c
		"11001110",	-- 0x3e0d
		"00111100",	-- 0x3e0e
		"00000001",	-- 0x3e0f
		"11001101",	-- 0x3e10
		"10001101",	-- 0x3e11
		"00000011",	-- 0x3e12
		"11111011",	-- 0x3e13
		"00011010",	-- 0x3e14
		"10110011",	-- 0x3e15
		"00000001",	-- 0x3e16
		"01010100",	-- 0x3e17
		"00110111",	-- 0x3e18
		"11010101",	-- 0x3e19
		"00001001",	-- 0x3e1a
		"01111001",	-- 0x3e1b
		"00011000",	-- 0x3e1c
		"10111001",	-- 0x3e1d
		"01000101",	-- 0x3e1e
		"00000100",	-- 0x3e1f
		"11001101",	-- 0x3e20
		"11110000",	-- 0x3e21
		"01000100",	-- 0x3e22
		"00001010",	-- 0x3e23
		"11111010",	-- 0x3e24
		"00000001",	-- 0x3e25
		"11011100",	-- 0x3e26
		"11000010",	-- 0x3e27
		"11111011",	-- 0x3e28
		"10110010",	-- 0x3e29
		"00000001",	-- 0x3e2a
		"11011100",	-- 0x3e2b
		"01000000",	-- 0x3e2c
		"00011011",	-- 0x3e2d
		"11111010",	-- 0x3e2e
		"00000001",	-- 0x3e2f
		"11011100",	-- 0x3e30
		"11000110",	-- 0x3e31
		"00000100",	-- 0x3e32
		"10110010",	-- 0x3e33
		"00000001",	-- 0x3e34
		"11011100",	-- 0x3e35
		"10000110",	-- 0x3e36
		"11111111",	-- 0x3e37
		"11111111",	-- 0x3e38
		"10111010",	-- 0x3e39
		"00000001",	-- 0x3e3a
		"01010010",	-- 0x3e3b
		"01110101",	-- 0x3e3c
		"01111100",	-- 0x3e3d
		"11111010",	-- 0x3e3e
		"00000001",	-- 0x3e3f
		"10001100",	-- 0x3e40
		"11000010",	-- 0x3e41
		"10111111",	-- 0x3e42
		"10110010",	-- 0x3e43
		"00000001",	-- 0x3e44
		"10001100",	-- 0x3e45
		"00000011",	-- 0x3e46
		"11111110",	-- 0x3e47
		"11100111",	-- 0x3e48
		"11111010",	-- 0x3e49
		"00000001",	-- 0x3e4a
		"10001100",	-- 0x3e4b
		"11001101",	-- 0x3e4c
		"00001101",	-- 0x3e4d
		"01000101",	-- 0x3e4e
		"00011010",	-- 0x3e4f
		"11001101",	-- 0x3e50
		"11111011",	-- 0x3e51
		"01000010",	-- 0x3e52
		"00011001",	-- 0x3e53
		"00110111",	-- 0x3e54
		"01011001",	-- 0x3e55
		"00001111",	-- 0x3e56
		"11001101",	-- 0x3e57
		"01001101",	-- 0x3e58
		"01000010",	-- 0x3e59
		"00010010",	-- 0x3e5a
		"11001101",	-- 0x3e5b
		"00110001",	-- 0x3e5c
		"01000010",	-- 0x3e5d
		"00000111",	-- 0x3e5e
		"11000010",	-- 0x3e5f
		"10111111",	-- 0x3e60
		"00110101",	-- 0x3e61
		"01010000",	-- 0x3e62
		"00000010",	-- 0x3e63
		"01110101",	-- 0x3e64
		"01111100",	-- 0x3e65
		"11000010",	-- 0x3e66
		"01111111",	-- 0x3e67
		"01000000",	-- 0x3e68
		"00011010",	-- 0x3e69
		"00110101",	-- 0x3e6a
		"01011001",	-- 0x3e6b
		"11111001",	-- 0x3e6c
		"11000110",	-- 0x3e6d
		"01000000",	-- 0x3e6e
		"11001110",	-- 0x3e6f
		"10000000",	-- 0x3e70
		"01000110",	-- 0x3e71
		"00000100",	-- 0x3e72
		"01110010",	-- 0x3e73
		"11011111",	-- 0x3e74
		"11000110",	-- 0x3e75
		"10000000",	-- 0x3e76
		"00110101",	-- 0x3e77
		"01010000",	-- 0x3e78
		"00000110",	-- 0x3e79
		"01111001",	-- 0x3e7a
		"00001111",	-- 0x3e7b
		"11011111",	-- 0x3e7c
		"01000101",	-- 0x3e7d
		"00000101",	-- 0x3e7e
		"10001100",	-- 0x3e7f
		"01110111",	-- 0x3e80
		"01111000",	-- 0x3e81
		"01110111",	-- 0x3e82
		"01111100",	-- 0x3e83
		"10110010",	-- 0x3e84
		"00000001",	-- 0x3e85
		"10001100",	-- 0x3e86
		"11001110",	-- 0x3e87
		"01000000",	-- 0x3e88
		"01000111",	-- 0x3e89
		"00000111",	-- 0x3e8a
		"10000110",	-- 0x3e8b
		"10100000",	-- 0x3e8c
		"01000010",	-- 0x3e8d
		"01110101",	-- 0x3e8e
		"10111101",	-- 0x3e8f
		"01000000",	-- 0x3e90
		"01010010",	-- 0x3e91
		"11001010",	-- 0x3e92
		"10101110",	-- 0x3e93
		"00110101",	-- 0x3e94
		"00010010",	-- 0x3e95
		"00000100",	-- 0x3e96
		"01110101",	-- 0x3e97
		"10111101",	-- 0x3e98
		"01000000",	-- 0x3e99
		"00111100",	-- 0x3e9a
		"00110111",	-- 0x3e9b
		"11010101",	-- 0x3e9c
		"00110100",	-- 0x3e9d
		"00111100",	-- 0x3e9e
		"00000001",	-- 0x3e9f
		"11000100",	-- 0x3ea0
		"11001010",	-- 0x3ea1
		"11110001",	-- 0x3ea2
		"00000011",	-- 0x3ea3
		"00000010",	-- 0x3ea4
		"10000000",	-- 0x3ea5
		"00000000",	-- 0x3ea6
		"00000100",	-- 0x3ea7
		"11110001",	-- 0x3ea8
		"00000011",	-- 0x3ea9
		"00000010",	-- 0x3eaa
		"10000000",	-- 0x3eab
		"00000000",	-- 0x3eac
		"00000100",	-- 0x3ead
		"01011000",	-- 0x3eae
		"01000111",	-- 0x3eaf
		"00000010",	-- 0x3eb0
		"11001011",	-- 0x3eb1
		"11111111",	-- 0x3eb2
		"11111010",	-- 0x3eb3
		"00000011",	-- 0x3eb4
		"00000010",	-- 0x3eb5
		"01110001",	-- 0x3eb6
		"10111101",	-- 0x3eb7
		"01000110",	-- 0x3eb8
		"00000110",	-- 0x3eb9
		"11000000",	-- 0x3eba
		"00000001",	-- 0x3ebb
		"01000100",	-- 0x3ebc
		"00000010",	-- 0x3ebd
		"11001010",	-- 0x3ebe
		"11111111",	-- 0x3ebf
		"00001011",	-- 0x3ec0
		"01000010",	-- 0x3ec1
		"00000001",	-- 0x3ec2
		"01011011",	-- 0x3ec3
		"10001111",	-- 0x3ec4
		"11000011",	-- 0x3ec5
		"11010101",	-- 0x3ec6
		"00100001",	-- 0x3ec7
		"10000010",	-- 0x3ec8
		"01101110",	-- 0x3ec9
		"10001110",	-- 0x3eca
		"00000011",	-- 0x3ecb
		"00000010",	-- 0x3ecc
		"00000001",	-- 0x3ecd
		"11010001",	-- 0x3ece
		"10011000",	-- 0x3ecf
		"01111110",	-- 0x3ed0
		"10001100",	-- 0x3ed1
		"01110101",	-- 0x3ed2
		"10111101",	-- 0x3ed3
		"11111010",	-- 0x3ed4
		"00000011",	-- 0x3ed5
		"00000010",	-- 0x3ed6
		"01010011",	-- 0x3ed7
		"00000100",	-- 0x3ed8
		"00000100",	-- 0x3ed9
		"01101000",	-- 0x3eda
		"00111100",	-- 0x3edb
		"00101110",	-- 0x3edc
		"10101000",	-- 0x3edd
		"00000000",	-- 0x3ede
		"01111110",	-- 0x3edf
		"01000100",	-- 0x3ee0
		"00000010",	-- 0x3ee1
		"01010010",	-- 0x3ee2
		"01010011",	-- 0x3ee3
		"10111010",	-- 0x3ee4
		"00000001",	-- 0x3ee5
		"01010010",	-- 0x3ee6
		"00000011",	-- 0x3ee7
		"11111011",	-- 0x3ee8
		"00011010",	-- 0x3ee9
		"10001111",	-- 0x3eea
		"11000011",	-- 0x3eeb
		"11001001",	-- 0x3eec
		"00100001",	-- 0x3eed
		"10001110",	-- 0x3eee
		"11111010",	-- 0x3eef
		"00000001",	-- 0x3ef0
		"10001100",	-- 0x3ef1
		"01000100",	-- 0x3ef2
		"00011001",	-- 0x3ef3
		"11001110",	-- 0x3ef4
		"00000100",	-- 0x3ef5
		"01000110",	-- 0x3ef6
		"00000100",	-- 0x3ef7
		"11000110",	-- 0x3ef8
		"00000100",	-- 0x3ef9
		"01110010",	-- 0x3efa
		"11011111",	-- 0x3efb
		"00110101",	-- 0x3efc
		"01010000",	-- 0x3efd
		"00000110",	-- 0x3efe
		"01111001",	-- 0x3eff
		"00001111",	-- 0x3f00
		"11011111",	-- 0x3f01
		"01000101",	-- 0x3f02
		"00000101",	-- 0x3f03
		"10001100",	-- 0x3f04
		"01110111",	-- 0x3f05
		"01111000",	-- 0x3f06
		"01110111",	-- 0x3f07
		"10011011",	-- 0x3f08
		"11001011",	-- 0x3f09
		"01111001",	-- 0x3f0a
		"01000000",	-- 0x3f0b
		"00000111",	-- 0x3f0c
		"00110101",	-- 0x3f0d
		"01010000",	-- 0x3f0e
		"00000010",	-- 0x3f0f
		"01110101",	-- 0x3f10
		"10011011",	-- 0x3f11
		"11000010",	-- 0x3f12
		"11111011",	-- 0x3f13
		"10110010",	-- 0x3f14
		"00000001",	-- 0x3f15
		"10001100",	-- 0x3f16
		"11001001",	-- 0x3f17
		"11111111",	-- 0x3f18
		"10010011",	-- 0x3f19
		"01010100",	-- 0x3f1a
		"10110011",	-- 0x3f1b
		"00000010",	-- 0x3f1c
		"00001010",	-- 0x3f1d
		"00000011",	-- 0x3f1e
		"11111011",	-- 0x3f1f
		"00011010",	-- 0x3f20
		"10001111",	-- 0x3f21
		"11000011",	-- 0x3f22
		"11001011",	-- 0x3f23
		"00100001",	-- 0x3f24
		"10001100",	-- 0x3f25
		"11111010",	-- 0x3f26
		"00000001",	-- 0x3f27
		"10001101",	-- 0x3f28
		"01000100",	-- 0x3f29
		"00011001",	-- 0x3f2a
		"11001110",	-- 0x3f2b
		"00000001",	-- 0x3f2c
		"01000110",	-- 0x3f2d
		"00000100",	-- 0x3f2e
		"11000110",	-- 0x3f2f
		"00000001",	-- 0x3f30
		"01110010",	-- 0x3f31
		"11011111",	-- 0x3f32
		"00110101",	-- 0x3f33
		"01010000",	-- 0x3f34
		"00000110",	-- 0x3f35
		"01111001",	-- 0x3f36
		"00001111",	-- 0x3f37
		"11011111",	-- 0x3f38
		"01000101",	-- 0x3f39
		"00000101",	-- 0x3f3a
		"10001100",	-- 0x3f3b
		"01110111",	-- 0x3f3c
		"01111000",	-- 0x3f3d
		"01110111",	-- 0x3f3e
		"10011100",	-- 0x3f3f
		"11001011",	-- 0x3f40
		"01111001",	-- 0x3f41
		"01000000",	-- 0x3f42
		"00000111",	-- 0x3f43
		"00110101",	-- 0x3f44
		"01010000",	-- 0x3f45
		"00000010",	-- 0x3f46
		"01110101",	-- 0x3f47
		"10011100",	-- 0x3f48
		"11000010",	-- 0x3f49
		"11111110",	-- 0x3f4a
		"10110010",	-- 0x3f4b
		"00000001",	-- 0x3f4c
		"10001101",	-- 0x3f4d
		"11001001",	-- 0x3f4e
		"11111111",	-- 0x3f4f
		"10010011",	-- 0x3f50
		"01010101",	-- 0x3f51
		"10110011",	-- 0x3f52
		"00000010",	-- 0x3f53
		"00001011",	-- 0x3f54
		"00000011",	-- 0x3f55
		"11111011",	-- 0x3f56
		"00011010",	-- 0x3f57
		"10010011",	-- 0x3f58
		"01010110",	-- 0x3f59
		"10110011",	-- 0x3f5a
		"00000010",	-- 0x3f5b
		"00001100",	-- 0x3f5c
		"00110111",	-- 0x3f5d
		"10101010",	-- 0x3f5e
		"00001010",	-- 0x3f5f
		"11001101",	-- 0x3f60
		"01010011",	-- 0x3f61
		"01000101",	-- 0x3f62
		"00000110",	-- 0x3f63
		"01110001",	-- 0x3f64
		"11010100",	-- 0x3f65
		"01000111",	-- 0x3f66
		"00000010",	-- 0x3f67
		"01110111",	-- 0x3f68
		"01000110",	-- 0x3f69
		"11011011",	-- 0x3f6a
		"01010110",	-- 0x3f6b
		"10001111",	-- 0x3f6c
		"11000001",	-- 0x3f6d
		"01000000",	-- 0x3f6e
		"00000001",	-- 0x3f6f
		"11000100",	-- 0x3f70
		"01000100",	-- 0x3f71
		"00000001",	-- 0x3f72
		"11000100",	-- 0x3f73
		"11001010",	-- 0x3f74
		"10111010",	-- 0x3f75
		"00000001",	-- 0x3f76
		"00011010",	-- 0x3f77
		"00000011",	-- 0x3f78
		"11111011",	-- 0x3f79
		"00011010",	-- 0x3f7a
		"10001111",	-- 0x3f7b
		"11000011",	-- 0x3f7c
		"11001101",	-- 0x3f7d
		"00100001",	-- 0x3f7e
		"10001010",	-- 0x3f7f
		"11111010",	-- 0x3f80
		"00000001",	-- 0x3f81
		"10001100",	-- 0x3f82
		"01000100",	-- 0x3f83
		"00011010",	-- 0x3f84
		"11001110",	-- 0x3f85
		"00000010",	-- 0x3f86
		"01000110",	-- 0x3f87
		"00000100",	-- 0x3f88
		"11000110",	-- 0x3f89
		"00000010",	-- 0x3f8a
		"01110010",	-- 0x3f8b
		"11011111",	-- 0x3f8c
		"00110101",	-- 0x3f8d
		"01010000",	-- 0x3f8e
		"00000110",	-- 0x3f8f
		"01111001",	-- 0x3f90
		"00001111",	-- 0x3f91
		"11011111",	-- 0x3f92
		"01000101",	-- 0x3f93
		"00000101",	-- 0x3f94
		"10001100",	-- 0x3f95
		"01110111",	-- 0x3f96
		"01111000",	-- 0x3f97
		"01110111",	-- 0x3f98
		"01111011",	-- 0x3f99
		"10001110",	-- 0x3f9a
		"00011011",	-- 0x3f9b
		"00000000",	-- 0x3f9c
		"01000000",	-- 0x3f9d
		"00000111",	-- 0x3f9e
		"00110101",	-- 0x3f9f
		"01010000",	-- 0x3fa0
		"00000010",	-- 0x3fa1
		"01110101",	-- 0x3fa2
		"01111011",	-- 0x3fa3
		"11000010",	-- 0x3fa4
		"11111101",	-- 0x3fa5
		"10110010",	-- 0x3fa6
		"00000001",	-- 0x3fa7
		"10001100",	-- 0x3fa8
		"00111100",	-- 0x3fa9
		"11001000",	-- 0x3faa
		"11111111",	-- 0x3fab
		"11001001",	-- 0x3fac
		"11111111",	-- 0x3fad
		"11000011",	-- 0x3fae
		"11000000",	-- 0x3faf
		"10011010",	-- 0x3fb0
		"01010111",	-- 0x3fb1
		"10111010",	-- 0x3fb2
		"00000010",	-- 0x3fb3
		"00000100",	-- 0x3fb4
		"00000011",	-- 0x3fb5
		"11111011",	-- 0x3fb6
		"00011010",	-- 0x3fb7
		"10110011",	-- 0x3fb8
		"00000001",	-- 0x3fb9
		"00000010",	-- 0x3fba
		"00000011",	-- 0x3fbb
		"11111011",	-- 0x3fbc
		"00011010",	-- 0x3fbd
		"10110011",	-- 0x3fbe
		"00000001",	-- 0x3fbf
		"11001011",	-- 0x3fc0
		"00000011",	-- 0x3fc1
		"11111011",	-- 0x3fc2
		"00011010",	-- 0x3fc3
		"10110011",	-- 0x3fc4
		"00000001",	-- 0x3fc5
		"11001100",	-- 0x3fc6
		"00000011",	-- 0x3fc7
		"11111011",	-- 0x3fc8
		"00011010",	-- 0x3fc9
		"10110011",	-- 0x3fca
		"00000001",	-- 0x3fcb
		"11001101",	-- 0x3fcc
		"00000011",	-- 0x3fcd
		"11111011",	-- 0x3fce
		"00011010",	-- 0x3fcf
		"10110011",	-- 0x3fd0
		"00000001",	-- 0x3fd1
		"11001110",	-- 0x3fd2
		"00000011",	-- 0x3fd3
		"11111011",	-- 0x3fd4
		"00011010",	-- 0x3fd5
		"00000011",	-- 0x3fd6
		"11111011",	-- 0x3fd7
		"00011010",	-- 0x3fd8
		"01011111",	-- 0x3fd9
		"01011111",	-- 0x3fda
		"11000100",	-- 0x3fdb
		"10000010",	-- 0x3fdc
		"10001000",	-- 0x3fdd
		"11111000",	-- 0x3fde
		"11110100",	-- 0x3fdf
		"11111010",	-- 0x3fe0
		"00001000",	-- 0x3fe1
		"11000000",	-- 0x3fe2
		"00000011",	-- 0x3fe3
		"11000000",	-- 0x3fe4
		"00000011",	-- 0x3fe5
		"11111001",	-- 0x3fe6
		"11000001",	-- 0x3fe7
		"11000000",	-- 0x3fe8
		"00000011",	-- 0x3fe9
		"11111001",	-- 0x3fea
		"10101100",	-- 0x3feb
		"11000000",	-- 0x3fec
		"00000011",	-- 0x3fed
		"11000000",	-- 0x3fee
		"00000011",	-- 0x3fef
		"11110110",	-- 0x3ff0
		"11110010",	-- 0x3ff1
		"11000000",	-- 0x3ff2
		"00000011",	-- 0x3ff3
		"11000000",	-- 0x3ff4
		"00000011",	-- 0x3ff5
		"11110111",	-- 0x3ff6
		"10011010",	-- 0x3ff7
		"11000000",	-- 0x3ff8
		"00000011",	-- 0x3ff9
		"11101111",	-- 0x3ffa
		"10110001",	-- 0x3ffb
		"11000000",	-- 0x3ffc
		"00000011",	-- 0x3ffd
		"11000110",	-- 0x3ffe
		"00000011");	-- 0x3fff
begin
	d <= rom(to_integer(unsigned(a))) when ce_n = '0' and oe_n = '0' else (others => 'Z');
end;
